H   �0�ŀ�@                        �5Gܞ$@                        rdB �G@H         0   �         `   �v�<w�<�v�<'w�<w�<�v�<w�<w�<�v�<,w�< w�<�v�<�v�<�v�< w�<,w�<�v�<w�<w�<�v�<w�<'w�<�v�<w�<`   `   w�<Aw�<w�<
w�<-w�<w�<w�<�v�<�v�<�v�<-w�<1w�<�v�<1w�<-w�<�v�<�v�<�v�<w�<w�<-w�<
w�<w�<Aw�<`   `   �v�<
w�<�v�<�v�<w�<�v�<w�<w�<w�<�v�<&w�<Yw�<�v�<Yw�<&w�<�v�<w�<w�<w�<�v�<w�<�v�<�v�<
w�<`   `   �v�<�v�<2w�<w�<w�<�v�<w�<	w�<w�<#w�<�v�<w�<�v�<w�<�v�<#w�<w�<	w�<w�<�v�<w�<w�<2w�<�v�<`   `   Aw�<w�<4w�<w�< w�<w�<$w�<�v�<�v�<3w�<�v�<(w�<w�<(w�<�v�<3w�<�v�<�v�<$w�<w�< w�<w�<4w�<w�<`   `   2w�<�v�<�v�<�v�<�v�<w�<w�<�v�<w�<#w�<�v�<w�<�v�<w�<�v�<#w�<w�<�v�<w�<w�<�v�<�v�<�v�<�v�<`   `   w�<+w�<w�<w�<$w�<w�<	w�<�v�<Aw�<�v�<�v�<w�<�v�<w�<�v�<�v�<Aw�<�v�<	w�<w�<$w�<w�<w�<+w�<`   `   w�<-w�<=w�<?w�<�v�<�v�<,w�<w�<w�<�v�<�v�<!w�<*w�<!w�<�v�<�v�<w�<w�<,w�<�v�<�v�<?w�<=w�<-w�<`   `   Iw�<w�<w�<&w�<�v�<�v�<w�<�v�<�v�<w�<w�<
w�<w�<
w�<w�<w�<�v�<�v�<w�<�v�<�v�<&w�<w�<w�<`   `   Ow�<�v�<w�< w�<w�<#w�<w�<#w�<w�<&w�<�v�<w�<(w�<w�<�v�<&w�<w�<#w�<w�<#w�<w�< w�<w�<�v�<`   `   �v�<�v�<0w�<�v�<.w�<&w�<7w�<@w�<�v�<w�<�v�<w�<�v�<w�<�v�<w�<�v�<@w�<7w�<&w�<.w�<�v�<0w�<�v�<`   `   6w�<w�<Pw�<w�<!w�<�v�<�v�<w�<�v�< w�<w�<w�<�v�<w�<w�< w�<�v�<w�<�v�<�v�<!w�<w�<Pw�<w�<`   `   w�<�v�<!w�<�v�<w�<"w�<�v�<w�<6w�<"w�<�v�<w�<�v�<w�<�v�<"w�<6w�<w�<�v�<"w�<w�<�v�<!w�<�v�<`   `   w�<�v�<.w�<�v�<�v�<Xw�<�v�<w�<+w�<w�<�v�<#w�<Ww�<#w�<�v�<w�<+w�<w�<�v�<Xw�<�v�<�v�<.w�<�v�<`   `   �w�<-w�<&w�<w�<�v�<w�<�v�<#w�<w�<w�<0w�<�v�<
w�<�v�<0w�<w�<w�<#w�<�v�<w�<�v�<w�<&w�<-w�<`   `   :w�<�v�<�v�<-w�<w�<w�<(w�<Mw�<w�<�v�<w�<�v�<�v�<�v�<w�<�v�<w�<Mw�<(w�<w�<w�<-w�<�v�<�v�<`   `   �v�<%w�<w�<w�<!w�<*w�<w�<�v�<�v�<�v�<w�<"w�<&w�<"w�<w�<�v�<�v�<�v�<w�<*w�<!w�<w�<w�<%w�<`   `   �v�<~w�<Dw�<�v�<w�<w�<w�<w�<*w�<'w�<w�<w�<w�<w�<w�<'w�<*w�<w�<w�<w�<w�<�v�<Dw�<~w�<`   `   �v�<+w�<�v�<�v�<"w�<�v�<w�<)w�<Ww�<w�<�v�<w�<w�<w�<�v�<w�<Ww�<)w�<w�<�v�<"w�<�v�<�v�<+w�<`   `   	w�<w�<�v�<#w�<w�<w�<!w�<�v�<+w�<�v�<�v�<.w�<�v�<.w�<�v�<�v�<+w�<�v�<!w�<w�<w�<#w�<�v�<w�<`   `   w�<"w�<w�<*w�<�v�<&w�<Hw�<w�<0w�<�v�<w�<w�<�v�<w�<w�<�v�<0w�<w�<Hw�<&w�<�v�<*w�<w�<"w�<`   `   �v�<�v�<w�< w�<w�<w�<w�<w�<#w�<w�<w�<w�<�v�<w�<w�<w�<#w�<w�<w�<w�<w�< w�<w�<�v�<`   `   ;w�<w�<w�<w�<w�<w�<w�<"w�<w�<'w�<�v�<w�<Ew�<w�<�v�<'w�<w�<"w�<w�<w�<w�<w�<w�<w�<`   `   gw�<�v�<3w�<w�<�v�<Lw�<8w�<�v�<�v�<w�<�v�<w�<w�<w�<�v�<w�<�v�<�v�<8w�<Lw�<�v�<w�<3w�<�v�<`   `   �v�<�v�< w�<,w�<�v�<w�<w�<�v�<w�<'w�<�v�<w�<�v�<w�<�v�<'w�<w�<�v�<w�<w�<�v�<,w�< w�<�v�<`   `   �v�<1w�<-w�<�v�<�v�<�v�<w�<w�<-w�<
w�<w�<Aw�<w�<Aw�<w�<
w�<-w�<w�<w�<�v�<�v�<�v�<-w�<1w�<`   `   �v�<Yw�<&w�<�v�<w�<w�<w�<�v�<w�<�v�<�v�<
w�<�v�<
w�<�v�<�v�<w�<�v�<w�<w�<w�<�v�<&w�<Yw�<`   `   �v�<w�<�v�<#w�<w�<	w�<w�<�v�<w�<w�<2w�<�v�<�v�<�v�<2w�<w�<w�<�v�<w�<	w�<w�<#w�<�v�<w�<`   `   w�<(w�<�v�<3w�<�v�<�v�<$w�<w�< w�<w�<4w�<w�<Aw�<w�<4w�<w�< w�<w�<$w�<�v�<�v�<3w�<�v�<(w�<`   `   �v�<w�<�v�<#w�<w�<�v�<w�<w�<�v�<�v�<�v�<�v�<2w�<�v�<�v�<�v�<�v�<w�<w�<�v�<w�<#w�<�v�<w�<`   `   �v�<w�<�v�<�v�<Aw�<�v�<	w�<w�<$w�<w�<w�<+w�<w�<+w�<w�<w�<$w�<w�<	w�<�v�<Aw�<�v�<�v�<w�<`   `   *w�<!w�<�v�<�v�<w�<w�<,w�<�v�<�v�<?w�<=w�<-w�<w�<-w�<=w�<?w�<�v�<�v�<,w�<w�<w�<�v�<�v�<!w�<`   `   w�<
w�<w�<w�<�v�<�v�<w�<�v�<�v�<&w�<w�<w�<Iw�<w�<w�<&w�<�v�<�v�<w�<�v�<�v�<w�<w�<
w�<`   `   (w�<w�<�v�<&w�<w�<#w�<w�<#w�<w�< w�<w�<�v�<Ow�<�v�<w�< w�<w�<#w�<w�<#w�<w�<&w�<�v�<w�<`   `   �v�<w�<�v�<w�<�v�<@w�<7w�<&w�<.w�<�v�<0w�<�v�<�v�<�v�<0w�<�v�<.w�<&w�<7w�<@w�<�v�<w�<�v�<w�<`   `   �v�<w�<w�< w�<�v�<w�<�v�<�v�<!w�<w�<Pw�<w�<6w�<w�<Pw�<w�<!w�<�v�<�v�<w�<�v�< w�<w�<w�<`   `   �v�<w�<�v�<"w�<6w�<w�<�v�<"w�<w�<�v�<!w�<�v�<w�<�v�<!w�<�v�<w�<"w�<�v�<w�<6w�<"w�<�v�<w�<`   `   Ww�<#w�<�v�<w�<+w�<w�<�v�<Xw�<�v�<�v�<.w�<�v�<w�<�v�<.w�<�v�<�v�<Xw�<�v�<w�<+w�<w�<�v�<#w�<`   `   
w�<�v�<0w�<w�<w�<#w�<�v�<w�<�v�<w�<&w�<-w�<�w�<-w�<&w�<w�<�v�<w�<�v�<#w�<w�<w�<0w�<�v�<`   `   �v�<�v�<w�<�v�<w�<Mw�<(w�<w�<w�<-w�<�v�<�v�<:w�<�v�<�v�<-w�<w�<w�<(w�<Mw�<w�<�v�<w�<�v�<`   `   &w�<"w�<w�<�v�<�v�<�v�<w�<*w�<!w�<w�<w�<%w�<�v�<%w�<w�<w�<!w�<*w�<w�<�v�<�v�<�v�<w�<"w�<`   `   w�<w�<w�<'w�<*w�<w�<w�<w�<w�<�v�<Dw�<~w�<�v�<~w�<Dw�<�v�<w�<w�<w�<w�<*w�<'w�<w�<w�<`   `   w�<w�<�v�<w�<Ww�<)w�<w�<�v�<"w�<�v�<�v�<+w�<�v�<+w�<�v�<�v�<"w�<�v�<w�<)w�<Ww�<w�<�v�<w�<`   `   �v�<.w�<�v�<�v�<+w�<�v�<!w�<w�<w�<#w�<�v�<w�<	w�<w�<�v�<#w�<w�<w�<!w�<�v�<+w�<�v�<�v�<.w�<`   `   �v�<w�<w�<�v�<0w�<w�<Hw�<&w�<�v�<*w�<w�<"w�<w�<"w�<w�<*w�<�v�<&w�<Hw�<w�<0w�<�v�<w�<w�<`   `   �v�<w�<w�<w�<#w�<w�<w�<w�<w�< w�<w�<�v�<�v�<�v�<w�< w�<w�<w�<w�<w�<#w�<w�<w�<w�<`   `   Ew�<w�<�v�<'w�<w�<"w�<w�<w�<w�<w�<w�<w�<;w�<w�<w�<w�<w�<w�<w�<"w�<w�<'w�<�v�<w�<`   `   w�<w�<�v�<w�<�v�<�v�<8w�<Lw�<�v�<w�<3w�<�v�<gw�<�v�<3w�<w�<�v�<Lw�<8w�<�v�<�v�<w�<�v�<w�<`   `   ow�<{w�<`w�<7w�<^w�<�w�<bw�<Tw�<�w�<Yw�<`w�<�w�<�w�<�w�<`w�<Yw�<�w�<Tw�<bw�<�w�<^w�<7w�<`w�<{w�<`   `   bw�<Hw�<mw�<�w�<Nw�<�w�<�w�<Zw�<�w�<ww�<,w�<jw�<�w�<jw�<,w�<ww�<�w�<Zw�<�w�<�w�<Nw�<�w�<mw�<Hw�<`   `   �w�<ew�<�w�<�w�<vw�<fw�<�w�<iw�<gw�<�w�<?w�<9w�<mw�<9w�<?w�<�w�<gw�<iw�<�w�<fw�<vw�<�w�<�w�<ew�<`   `   �w�<^w�<Kw�<hw�<�w�<^w�<^w�<�w�<Nw�<xw�<rw�<dw�<�w�<dw�<rw�<xw�<Nw�<�w�<^w�<^w�<�w�<hw�<Kw�<^w�<`   `   �w�<^w�<Uw�<Uw�<�w�<Tw�<Sw�<�w�<ow�<\w�<mw�<hw�<�w�<hw�<mw�<\w�<ow�<�w�<Sw�<Tw�<�w�<Uw�<Uw�<^w�<`   `   Pw�<tw�<�w�<�w�<�w�<gw�<|w�<�w�<^w�<Uw�<w�<jw�<~w�<jw�<w�<Uw�<^w�<�w�<|w�<gw�<�w�<�w�<�w�<tw�<`   `   :w�<tw�<�w�<ew�<ww�<nw�<jw�<qw�<4w�<�w�<�w�<sw�<�w�<sw�<�w�<�w�<4w�<qw�<jw�<nw�<ww�<ew�<�w�<tw�<`   `   <w�<Yw�<4w�<$w�<ww�<�w�<\w�<nw�<]w�<�w�<�w�<Cw�<hw�<Cw�<�w�<�w�<]w�<nw�<\w�<�w�<ww�<$w�<4w�<Yw�<`   `   Gw�<Tw�<^w�<fw�<�w�<�w�<]w�<�w�<rw�<^w�<�w�<Xw�<]w�<Xw�<�w�<^w�<rw�<�w�<]w�<�w�<�w�<fw�<^w�<Tw�<`   `   mw�<~w�<�w�<�w�<lw�<Sw�<+w�<\w�<[w�<Vw�<�w�<}w�<Iw�<}w�<�w�<Vw�<[w�<\w�<+w�<Sw�<lw�<�w�<�w�<~w�<`   `   ]w�<iw�<lw�<Tw�<ew�<gw�<Ww�<Uw�<{w�<|w�<pw�<yw�<Yw�<yw�<pw�<|w�<{w�<Uw�<Ww�<gw�<ew�<Tw�<lw�<iw�<`   `   lw�<Sw�<0w�<Nw�<w�<�w�<�w�<mw�<~w�<mw�<Ow�<�w�<�w�<�w�<Ow�<mw�<~w�<mw�<�w�<�w�<w�<Nw�<0w�<Sw�<`   `   �w�<�w�<Jw�<qw�<ww�<Dw�<�w�<zw�<Qw�<\w�<ow�<�w�<nw�<�w�<ow�<\w�<Qw�<zw�<�w�<Dw�<ww�<qw�<Jw�<�w�<`   `   [w�<w�<_w�<~w�<�w�<0w�<}w�<�w�<8w�<nw�<�w�<Cw�<w�<Cw�<�w�<nw�<8w�<�w�<}w�<0w�<�w�<~w�<_w�<w�<`   `   �v�<Ww�<\w�<\w�<�w�<^w�<w�<bw�<9w�<tw�<`w�<mw�<�w�<mw�<`w�<tw�<9w�<bw�<w�<^w�<�w�<\w�<\w�<Ww�<`   `   Yw�<�w�<�w�<Vw�<hw�<hw�<{w�<Pw�<vw�<�w�<[w�<�w�<�w�<�w�<[w�<�w�<vw�<Pw�<{w�<hw�<hw�<Vw�<�w�<�w�<`   `   �w�<uw�<dw�<pw�<Ew�<?w�<aw�<gw�<�w�<�w�<nw�<nw�<Iw�<nw�<nw�<�w�<�w�<gw�<aw�<?w�<Ew�<pw�<dw�<uw�<`   `   vw�<w�<,w�<�w�<fw�<Gw�<kw�<zw�<Xw�<Uw�<yw�<Zw�<)w�<Zw�<yw�<Uw�<Xw�<zw�<kw�<Gw�<fw�<�w�<,w�<w�<`   `   �w�<Uw�<tw�<�w�<yw�<vw�<�w�<iw�<w�<Vw�<�w�<yw�<�w�<yw�<�w�<Vw�<w�<iw�<�w�<vw�<yw�<�w�<tw�<Uw�<`   `   �w�<cw�<�w�<�w�<Pw�<vw�<aw�<Vw�<bw�<�w�<�w�<Xw�<�w�<Xw�<�w�<�w�<bw�<Vw�<aw�<vw�<Pw�<�w�<�w�<cw�<`   `   _w�<^w�<Kw�<Aw�<]w�<tw�<Iw�<Ow�<sw�<�w�<Vw�<Yw�<�w�<Yw�<Vw�<�w�<sw�<Ow�<Iw�<tw�<]w�<Aw�<Kw�<^w�<`   `   �w�<�w�<Uw�<Gw�<�w�<ww�<Xw�<Sw�<4w�<Vw�<Tw�<`w�<�w�<`w�<Tw�<Vw�<4w�<Sw�<Xw�<ww�<�w�<Gw�<Uw�<�w�<`   `   <w�<pw�<ow�<Xw�<�w�<^w�<Rw�<uw�<Vw�<|w�<�w�<Rw�<2w�<Rw�<�w�<|w�<Vw�<uw�<Rw�<^w�<�w�<Xw�<ow�<pw�<`   `   #w�<_w�<|w�<Uw�<zw�<Lw�<Aw�<�w�<�w�<sw�<�w�<�w�<Qw�<�w�<�w�<sw�<�w�<�w�<Aw�<Lw�<zw�<Uw�<|w�<_w�<`   `   �w�<�w�<`w�<Yw�<�w�<Tw�<bw�<�w�<^w�<7w�<`w�<{w�<ow�<{w�<`w�<7w�<^w�<�w�<bw�<Tw�<�w�<Yw�<`w�<�w�<`   `   �w�<jw�<,w�<ww�<�w�<Zw�<�w�<�w�<Nw�<�w�<mw�<Hw�<bw�<Hw�<mw�<�w�<Nw�<�w�<�w�<Zw�<�w�<ww�<,w�<jw�<`   `   mw�<9w�<?w�<�w�<gw�<iw�<�w�<fw�<vw�<�w�<�w�<ew�<�w�<ew�<�w�<�w�<vw�<fw�<�w�<iw�<gw�<�w�<?w�<9w�<`   `   �w�<dw�<rw�<xw�<Nw�<�w�<^w�<^w�<�w�<hw�<Kw�<^w�<�w�<^w�<Kw�<hw�<�w�<^w�<^w�<�w�<Nw�<xw�<rw�<dw�<`   `   �w�<hw�<mw�<\w�<ow�<�w�<Sw�<Tw�<�w�<Uw�<Uw�<^w�<�w�<^w�<Uw�<Uw�<�w�<Tw�<Sw�<�w�<ow�<\w�<mw�<hw�<`   `   ~w�<jw�<w�<Uw�<^w�<�w�<|w�<gw�<�w�<�w�<�w�<tw�<Pw�<tw�<�w�<�w�<�w�<gw�<|w�<�w�<^w�<Uw�<w�<jw�<`   `   �w�<sw�<�w�<�w�<4w�<qw�<jw�<nw�<ww�<ew�<�w�<tw�<:w�<tw�<�w�<ew�<ww�<nw�<jw�<qw�<4w�<�w�<�w�<sw�<`   `   hw�<Cw�<�w�<�w�<]w�<nw�<\w�<�w�<ww�<$w�<4w�<Yw�<<w�<Yw�<4w�<$w�<ww�<�w�<\w�<nw�<]w�<�w�<�w�<Cw�<`   `   ]w�<Xw�<�w�<^w�<rw�<�w�<]w�<�w�<�w�<fw�<^w�<Tw�<Gw�<Tw�<^w�<fw�<�w�<�w�<]w�<�w�<rw�<^w�<�w�<Xw�<`   `   Iw�<}w�<�w�<Vw�<[w�<\w�<+w�<Sw�<lw�<�w�<�w�<~w�<mw�<~w�<�w�<�w�<lw�<Sw�<+w�<\w�<[w�<Vw�<�w�<}w�<`   `   Yw�<yw�<pw�<|w�<{w�<Uw�<Ww�<gw�<ew�<Tw�<lw�<iw�<]w�<iw�<lw�<Tw�<ew�<gw�<Ww�<Uw�<{w�<|w�<pw�<yw�<`   `   �w�<�w�<Ow�<mw�<~w�<mw�<�w�<�w�<w�<Nw�<0w�<Sw�<lw�<Sw�<0w�<Nw�<w�<�w�<�w�<mw�<~w�<mw�<Ow�<�w�<`   `   nw�<�w�<ow�<\w�<Qw�<zw�<�w�<Dw�<ww�<qw�<Jw�<�w�<�w�<�w�<Jw�<qw�<ww�<Dw�<�w�<zw�<Qw�<\w�<ow�<�w�<`   `   w�<Cw�<�w�<nw�<8w�<�w�<}w�<0w�<�w�<~w�<_w�<w�<[w�<w�<_w�<~w�<�w�<0w�<}w�<�w�<8w�<nw�<�w�<Cw�<`   `   �w�<mw�<`w�<tw�<9w�<bw�<w�<^w�<�w�<\w�<\w�<Ww�<�v�<Ww�<\w�<\w�<�w�<^w�<w�<bw�<9w�<tw�<`w�<mw�<`   `   �w�<�w�<[w�<�w�<vw�<Pw�<{w�<hw�<hw�<Vw�<�w�<�w�<Yw�<�w�<�w�<Vw�<hw�<hw�<{w�<Pw�<vw�<�w�<[w�<�w�<`   `   Iw�<nw�<nw�<�w�<�w�<gw�<aw�<?w�<Ew�<pw�<dw�<uw�<�w�<uw�<dw�<pw�<Ew�<?w�<aw�<gw�<�w�<�w�<nw�<nw�<`   `   )w�<Zw�<yw�<Uw�<Xw�<zw�<kw�<Gw�<fw�<�w�<,w�<w�<vw�<w�<,w�<�w�<fw�<Gw�<kw�<zw�<Xw�<Uw�<yw�<Zw�<`   `   �w�<yw�<�w�<Vw�<w�<iw�<�w�<vw�<yw�<�w�<tw�<Uw�<�w�<Uw�<tw�<�w�<yw�<vw�<�w�<iw�<w�<Vw�<�w�<yw�<`   `   �w�<Xw�<�w�<�w�<bw�<Vw�<aw�<vw�<Pw�<�w�<�w�<cw�<�w�<cw�<�w�<�w�<Pw�<vw�<aw�<Vw�<bw�<�w�<�w�<Xw�<`   `   �w�<Yw�<Vw�<�w�<sw�<Ow�<Iw�<tw�<]w�<Aw�<Kw�<^w�<_w�<^w�<Kw�<Aw�<]w�<tw�<Iw�<Ow�<sw�<�w�<Vw�<Yw�<`   `   �w�<`w�<Tw�<Vw�<4w�<Sw�<Xw�<ww�<�w�<Gw�<Uw�<�w�<�w�<�w�<Uw�<Gw�<�w�<ww�<Xw�<Sw�<4w�<Vw�<Tw�<`w�<`   `   2w�<Rw�<�w�<|w�<Vw�<uw�<Rw�<^w�<�w�<Xw�<ow�<pw�<<w�<pw�<ow�<Xw�<�w�<^w�<Rw�<uw�<Vw�<|w�<�w�<Rw�<`   `   Qw�<�w�<�w�<sw�<�w�<�w�<Aw�<Lw�<zw�<Uw�<|w�<_w�<#w�<_w�<|w�<Uw�<zw�<Lw�<Aw�<�w�<�w�<sw�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<x�<�w�< x�<�w�<x�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   $x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�< x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<`   `   �w�<�w�<�w�< x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�< x�<�w�<�w�<`   `   w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<x�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�< x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�< x�<�w�<�w�<`   `   �w�<�w�<�w�<x�<�w�<�w�<x�<	x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<	x�<x�<�w�<�w�<x�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<`   `   �w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<`   `    x�<�w�<x�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<x�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<$x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `    x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�< x�<�w�<�w�<�w�<�w�<�w�< x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�< x�<�w�<�w�<�w�<�w�<�w�< x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<	x�<x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<x�<	x�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   /x�<@x�<{x�<qx�<[x�<Hx�<nx�<Ux�<0x�<[x�<=x�<<x�<8x�<<x�<=x�<[x�<0x�<Ux�<nx�<Hx�<[x�<qx�<{x�<@x�<`   `   Zx�<qx�<Qx�<6x�<zx�<fx�<?x�<dx�<>x�<Bx�<`x�<Qx�<^x�<Qx�<`x�<Bx�<>x�<dx�<?x�<fx�<zx�<6x�<Qx�<qx�<`   `   6x�<dx�<'x�<)x�<ix�<Wx�<-x�<dx�<jx�<x�<2x�<Nx�<�x�<Nx�<2x�<x�<jx�<dx�<-x�<Wx�<ix�<)x�<'x�<dx�<`   `   $x�<ax�<Qx�<�x�<9x�<x�<ax�<kx�<�x�<x�<x�<,x�<,x�<,x�<x�<x�<�x�<kx�<ax�<x�<9x�<�x�<Qx�<ax�<`   `   Rx�<ex�<Cx�<�x�<>x�</x�<|x�<<x�<xx�<Ix�<Vx�<dx�<>x�<dx�<Vx�<Ix�<xx�<<x�<|x�</x�<>x�<�x�<Cx�<ex�<`   `   tx�<Zx�<x�<Sx�<Gx�<Sx�<dx�<&x�<lx�<Wx�<Wx�<�x�<ox�<�x�<Wx�<Wx�<lx�<&x�<dx�<Sx�<Gx�<Sx�<x�<Zx�<`   `   3x�<!x�<9x�<ax�<bx�<ox�<vx�<kx�<vx�<Gx�<Px�<`x�<$x�<`x�<Px�<Gx�<vx�<kx�<vx�<ox�<bx�<ax�<9x�<!x�<`   `   x�<x�<Wx�<ux�<^x�<Yx�<Yx�<Ax�<Jx�<Cx�<vx�<vx�<x�<vx�<vx�<Cx�<Jx�<Ax�<Yx�<Yx�<^x�<ux�<Wx�<x�<`   `   >x�<Qx�<Fx�<?x�<)x�<-x�<8x�<�w�<Kx�<qx�<Zx�<Jx�<x�<Jx�<Zx�<qx�<Kx�<�w�<8x�<-x�<)x�<?x�<Fx�<Qx�<`   `   ,x�<Ox�<.x�<]x�<`x�<Px�<^x�<(x�<Vx�<px�<=x�<$x�<Dx�<$x�<=x�<px�<Vx�<(x�<^x�<Px�<`x�<]x�<.x�<Ox�<`   `   Rx�<]x�<*x�<lx�<qx�<Lx�<Hx�<\x�<'x�<*x�<}x�<hx�<�x�<hx�<}x�<*x�<'x�<\x�<Hx�<Lx�<qx�<lx�<*x�<]x�<`   `   nx�<mx�<5x�<5x�<7x�<Qx�<0x�<�x�<Kx�<-x�<�x�<Kx�<qx�<Kx�<�x�<-x�<Kx�<�x�<0x�<Qx�<7x�<5x�<5x�<mx�<`   `   =x�<7x�<7x�<7x�<?x�<�x�<:x�<[x�<]x�<1x�<ax�<+x�<Tx�<+x�<ax�<1x�<]x�<[x�<:x�<�x�<?x�<7x�<7x�<7x�<`   `   lx�<+x�<1x�<Px�<8x�<�x�<Ex�<+x�<Gx�<x�<*x�<`x�<�x�<`x�<*x�<x�<Gx�<+x�<Ex�<�x�<8x�<Px�<1x�<+x�<`   `   �x�<Fx�<Rx�<qx�<+x�<Kx�<Lx�<Rx�<Xx�<%x�<Lx�<jx�<Fx�<jx�<Lx�<%x�<Xx�<Rx�<Lx�<Kx�<+x�<qx�<Rx�<Fx�<`   `   dx�<x�<@x�<Vx�<3x�<+x�<Lx�<wx�<Bx�<Ix�<�x�<lx�<0x�<lx�<�x�<Ix�<Bx�<wx�<Lx�<+x�<3x�<Vx�<@x�<x�<`   `   Sx�<9x�<Cx�<!x�<8x�<5x�<Ux�<zx�<'x�<Ex�<ax�<jx�<ox�<jx�<ax�<Ex�<'x�<zx�<Ux�<5x�<8x�<!x�<Cx�<9x�<`   `   Ex�<yx�<�x�<Bx�<Sx�<>x�<:x�<@x�<Fx�<gx�<1x�<5x�<7x�<5x�<1x�<gx�<Fx�<@x�<:x�<>x�<Sx�<Bx�<�x�<yx�<`   `   �w�<<x�<]x�<Kx�<px�<Dx�<Gx�<;x�<kx�<vx�<?x�<Fx�<x�<Fx�<?x�<vx�<kx�<;x�<Gx�<Dx�<px�<Kx�<]x�<<x�<`   `   ax�<Mx�<"x�<Qx�<�x�<Cx�<_x�<Jx�<:x�<,x�<Wx�<�x�<ax�<�x�<Wx�<,x�<:x�<Jx�<_x�<Cx�<�x�<Qx�<"x�<Mx�<`   `   �x�<mx�<?x�<Ox�<Tx�<Ex�<;x�<x�<x�<#x�<[x�<jx�< x�<jx�<[x�<#x�<x�<x�<;x�<Ex�<Tx�<Ox�<?x�<mx�<`   `   $x�<)x�<0x�<(x�<x�<fx�<;x�<x�<cx�<bx�<dx�<Bx�<x�<Bx�<dx�<bx�<cx�<x�<;x�<fx�<x�<(x�<0x�<)x�<`   `   dx�<Px�<0x�<_x�<9x�<ax�<Nx�<x�<fx�<Gx�<Nx�<qx�<�x�<qx�<Nx�<Gx�<fx�<x�<Nx�<ax�<9x�<_x�<0x�<Px�<`   `   �x�<kx�</x�<�x�<Px�<Fx�<ix�<.x�<Gx�<Ix�<Kx�<>x�<Wx�<>x�<Kx�<Ix�<Gx�<.x�<ix�<Fx�<Px�<�x�</x�<kx�<`   `   8x�<<x�<=x�<[x�<0x�<Ux�<nx�<Hx�<[x�<qx�<{x�<@x�</x�<@x�<{x�<qx�<[x�<Hx�<nx�<Ux�<0x�<[x�<=x�<<x�<`   `   ^x�<Qx�<`x�<Bx�<>x�<dx�<?x�<fx�<zx�<6x�<Qx�<qx�<Zx�<qx�<Qx�<6x�<zx�<fx�<?x�<dx�<>x�<Bx�<`x�<Qx�<`   `   �x�<Nx�<2x�<x�<jx�<dx�<-x�<Wx�<ix�<)x�<'x�<dx�<6x�<dx�<'x�<)x�<ix�<Wx�<-x�<dx�<jx�<x�<2x�<Nx�<`   `   ,x�<,x�<x�<x�<�x�<kx�<ax�<x�<9x�<�x�<Qx�<ax�<$x�<ax�<Qx�<�x�<9x�<x�<ax�<kx�<�x�<x�<x�<,x�<`   `   >x�<dx�<Vx�<Ix�<xx�<<x�<|x�</x�<>x�<�x�<Cx�<ex�<Rx�<ex�<Cx�<�x�<>x�</x�<|x�<<x�<xx�<Ix�<Vx�<dx�<`   `   ox�<�x�<Wx�<Wx�<lx�<&x�<dx�<Sx�<Gx�<Sx�<x�<Zx�<tx�<Zx�<x�<Sx�<Gx�<Sx�<dx�<&x�<lx�<Wx�<Wx�<�x�<`   `   $x�<`x�<Px�<Gx�<vx�<kx�<vx�<ox�<bx�<ax�<9x�<!x�<3x�<!x�<9x�<ax�<bx�<ox�<vx�<kx�<vx�<Gx�<Px�<`x�<`   `   x�<vx�<vx�<Cx�<Jx�<Ax�<Yx�<Yx�<^x�<ux�<Wx�<x�<x�<x�<Wx�<ux�<^x�<Yx�<Yx�<Ax�<Jx�<Cx�<vx�<vx�<`   `   x�<Jx�<Zx�<qx�<Kx�<�w�<8x�<-x�<)x�<?x�<Fx�<Qx�<>x�<Qx�<Fx�<?x�<)x�<-x�<8x�<�w�<Kx�<qx�<Zx�<Jx�<`   `   Dx�<$x�<=x�<px�<Vx�<(x�<^x�<Px�<`x�<]x�<.x�<Ox�<,x�<Ox�<.x�<]x�<`x�<Px�<^x�<(x�<Vx�<px�<=x�<$x�<`   `   �x�<hx�<}x�<*x�<'x�<\x�<Hx�<Lx�<qx�<lx�<*x�<]x�<Rx�<]x�<*x�<lx�<qx�<Lx�<Hx�<\x�<'x�<*x�<}x�<hx�<`   `   qx�<Kx�<�x�<-x�<Kx�<�x�<0x�<Qx�<7x�<5x�<5x�<mx�<nx�<mx�<5x�<5x�<7x�<Qx�<0x�<�x�<Kx�<-x�<�x�<Kx�<`   `   Tx�<+x�<ax�<1x�<]x�<[x�<:x�<�x�<?x�<7x�<7x�<7x�<=x�<7x�<7x�<7x�<?x�<�x�<:x�<[x�<]x�<1x�<ax�<+x�<`   `   �x�<`x�<*x�<x�<Gx�<+x�<Ex�<�x�<8x�<Px�<1x�<+x�<lx�<+x�<1x�<Px�<8x�<�x�<Ex�<+x�<Gx�<x�<*x�<`x�<`   `   Fx�<jx�<Lx�<%x�<Xx�<Rx�<Lx�<Kx�<+x�<qx�<Rx�<Fx�<�x�<Fx�<Rx�<qx�<+x�<Kx�<Lx�<Rx�<Xx�<%x�<Lx�<jx�<`   `   0x�<lx�<�x�<Ix�<Bx�<wx�<Lx�<+x�<3x�<Vx�<@x�<x�<dx�<x�<@x�<Vx�<3x�<+x�<Lx�<wx�<Bx�<Ix�<�x�<lx�<`   `   ox�<jx�<ax�<Ex�<'x�<zx�<Ux�<5x�<8x�<!x�<Cx�<9x�<Sx�<9x�<Cx�<!x�<8x�<5x�<Ux�<zx�<'x�<Ex�<ax�<jx�<`   `   7x�<5x�<1x�<gx�<Fx�<@x�<:x�<>x�<Sx�<Bx�<�x�<yx�<Ex�<yx�<�x�<Bx�<Sx�<>x�<:x�<@x�<Fx�<gx�<1x�<5x�<`   `   x�<Fx�<?x�<vx�<kx�<;x�<Gx�<Dx�<px�<Kx�<]x�<<x�<�w�<<x�<]x�<Kx�<px�<Dx�<Gx�<;x�<kx�<vx�<?x�<Fx�<`   `   ax�<�x�<Wx�<,x�<:x�<Jx�<_x�<Cx�<�x�<Qx�<"x�<Mx�<ax�<Mx�<"x�<Qx�<�x�<Cx�<_x�<Jx�<:x�<,x�<Wx�<�x�<`   `    x�<jx�<[x�<#x�<x�<x�<;x�<Ex�<Tx�<Ox�<?x�<mx�<�x�<mx�<?x�<Ox�<Tx�<Ex�<;x�<x�<x�<#x�<[x�<jx�<`   `   x�<Bx�<dx�<bx�<cx�<x�<;x�<fx�<x�<(x�<0x�<)x�<$x�<)x�<0x�<(x�<x�<fx�<;x�<x�<cx�<bx�<dx�<Bx�<`   `   �x�<qx�<Nx�<Gx�<fx�<x�<Nx�<ax�<9x�<_x�<0x�<Px�<dx�<Px�<0x�<_x�<9x�<ax�<Nx�<x�<fx�<Gx�<Nx�<qx�<`   `   Wx�<>x�<Kx�<Ix�<Gx�<.x�<ix�<Fx�<Px�<�x�</x�<kx�<�x�<kx�</x�<�x�<Px�<Fx�<ix�<.x�<Gx�<Ix�<Kx�<>x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<y�<*y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<*y�<y�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<y�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<y�<`   `   }x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�< y�<�x�<y�<y�<�x�<�x�<�x�<�x�<�x�<y�<y�<�x�< y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�< y�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�< y�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�< y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�< y�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<*y�<y�<�x�<y�<*y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<y�<�x�<y�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<}x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   y�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<y�<y�<�x�< y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�< y�<�x�<y�<y�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�< y�<�x�<�x�<�x�< y�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�< y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�< y�<�x�<�x�<�x�<�x�<`   `   �y�<xy�<Iy�<�y�<�y�<Wy�<]y�<|y�<my�<my�<�y�<�y�<py�<�y�<�y�<my�<my�<|y�<]y�<Wy�<�y�<�y�<Iy�<xy�<`   `   qy�<Vy�<ky�<�y�<my�<Hy�<hy�<my�<?y�<Dy�<Wy�<[y�<By�<[y�<Wy�<Dy�<?y�<my�<hy�<Hy�<my�<�y�<ky�<Vy�<`   `   Ry�<@y�<uy�<my�<;y�<gy�<�y�<�y�<]y�<By�<\y�<Xy�<8y�<Xy�<\y�<By�<]y�<�y�<�y�<gy�<;y�<my�<uy�<@y�<`   `   �y�<wy�<�y�<Dy�<Hy�<~y�<By�<dy�<|y�<Zy�<Sy�<sy�<�y�<sy�<Sy�<Zy�<|y�<dy�<By�<~y�<Hy�<Dy�<�y�<wy�<`   `   ^y�<xy�<�y�<Fy�<ny�<}y�<4y�<�y�<�y�<fy�<=y�<;y�<ry�<;y�<=y�<fy�<�y�<�y�<4y�<}y�<ny�<Fy�<�y�<xy�<`   `   Hy�<9y�<ry�<Uy�<|y�<y�<ey�<�y�<hy�<�y�<�y�<`y�<xy�<`y�<�y�<�y�<hy�<�y�<ey�<y�<|y�<Uy�<ry�<9y�<`   `   �y�<y�<Ky�<ay�<ny�<�y�<uy�<ly�<Zy�<�y�<gy�<{y�<�y�<{y�<gy�<�y�<Zy�<ly�<uy�<�y�<ny�<ay�<Ky�<y�<`   `   �y�<2y�<�y�<�y�<iy�<^y�<^y�<_y�<oy�<�y�<.y�<Ay�<qy�<Ay�<.y�<�y�<oy�<_y�<^y�<^y�<iy�<�y�<�y�<2y�<`   `   Fy�<+y�<xy�<�y�<zy�<7y�<@y�<]y�<9y�<uy�<dy�<Yy�<Iy�<Yy�<dy�<uy�<9y�<]y�<@y�<7y�<zy�<�y�<xy�<+y�<`   `   py�<>y�<>y�<<y�<cy�<cy�<ay�<ay�<5y�<Oy�<�y�<�y�<]y�<�y�<�y�<Oy�<5y�<ay�<ay�<cy�<cy�<<y�<>y�<>y�<`   `   �y�<qy�<ty�<by�<Ny�<�y�<|y�<Jy�<�y�<�y�<my�<�y�<:y�<�y�<my�<�y�<�y�<Jy�<|y�<�y�<Ny�<by�<ty�<qy�<`   `   ay�<Ky�<ry�<�y�<my�<}y�<�y�<*y�<ny�<zy�<By�<}y�<Sy�<}y�<By�<zy�<ny�<*y�<�y�<}y�<my�<�y�<ry�<Ky�<`   `   <y�<Vy�<Ay�<7y�<vy�<Gy�<�y�<My�<<y�<Sy�<6y�<�y�<�y�<�y�<6y�<Sy�<<y�<My�<�y�<Gy�<vy�<7y�<Ay�<Vy�<`   `   \y�<�y�<Vy�<-y�<�y�<Fy�<�y�<{y�<Wy�<^y�<Ey�<�y�<Xy�<�y�<Ey�<^y�<Wy�<{y�<�y�<Fy�<�y�<-y�<Vy�<�y�<`   `   py�<~y�<Ey�<*y�<vy�<`y�<vy�<|y�<ay�<Gy�<Zy�<�y�<jy�<�y�<Zy�<Gy�<ay�<|y�<vy�<`y�<vy�<*y�<Ey�<~y�<`   `   ny�<{y�<Sy�<5y�<7y�<Ry�<_y�<fy�<Wy�<9y�<cy�<�y�<�y�<�y�<cy�<9y�<Wy�<fy�<_y�<Ry�<7y�<5y�<Sy�<{y�<`   `   2y�<ny�<�y�<y�<Gy�<jy�<cy�<^y�<jy�<_y�<|y�<;y�<Dy�<;y�<|y�<_y�<jy�<^y�<cy�<jy�<Gy�<y�<�y�<ny�<`   `   Ry�<py�<]y�<py�<Gy�<ry�<\y�<oy�<�y�<Ty�<�y�<{y�<�y�<{y�<�y�<Ty�<�y�<oy�<\y�<ry�<Gy�<py�<]y�<py�<`   `   y�<�y�<gy�<Ny�<Sy�<~y�<?y�<ky�<�y�<7y�<Yy�<fy�<yy�<fy�<Yy�<7y�<�y�<ky�<?y�<~y�<Sy�<Ny�<gy�<�y�<`   `   /y�<ky�<�y�<My�<xy�<�y�<6y�<:y�<Oy�<`y�<`y�<+y�<-y�<+y�<`y�<`y�<Oy�<:y�<6y�<�y�<xy�<My�<�y�<ky�<`   `   @y�<,y�<[y�<My�<uy�<ly�<Ly�<^y�<y�<py�<�y�<uy�<�y�<uy�<�y�<py�<y�<^y�<Ly�<ly�<uy�<My�<[y�<,y�<`   `   �y�<Gy�<Ly�<my�<iy�<2y�<Hy�<�y�<#y�<^y�<~y�<|y�<�y�<|y�<~y�<^y�<#y�<�y�<Hy�<2y�<iy�<my�<Ly�<Gy�<`   `   �y�<Xy�<[y�<Dy�<Qy�<ay�<Ny�<=y�<-y�<y�<vy�<Ty�<Ey�<Ty�<vy�<y�<-y�<=y�<Ny�<ay�<Qy�<Dy�<[y�<Xy�<`   `   By�<cy�<ty�<>y�<ly�<�y�<�y�<By�<ey�<�y�<[y�<_y�<xy�<_y�<[y�<�y�<ey�<By�<�y�<�y�<ly�<>y�<ty�<cy�<`   `   py�<�y�<�y�<my�<my�<|y�<]y�<Wy�<�y�<�y�<Iy�<xy�<�y�<xy�<Iy�<�y�<�y�<Wy�<]y�<|y�<my�<my�<�y�<�y�<`   `   By�<[y�<Wy�<Dy�<?y�<my�<hy�<Hy�<my�<�y�<ky�<Vy�<qy�<Vy�<ky�<�y�<my�<Hy�<hy�<my�<?y�<Dy�<Wy�<[y�<`   `   8y�<Xy�<\y�<By�<]y�<�y�<�y�<gy�<;y�<my�<uy�<@y�<Ry�<@y�<uy�<my�<;y�<gy�<�y�<�y�<]y�<By�<\y�<Xy�<`   `   �y�<sy�<Sy�<Zy�<|y�<dy�<By�<~y�<Hy�<Dy�<�y�<wy�<�y�<wy�<�y�<Dy�<Hy�<~y�<By�<dy�<|y�<Zy�<Sy�<sy�<`   `   ry�<;y�<=y�<fy�<�y�<�y�<4y�<}y�<ny�<Fy�<�y�<xy�<^y�<xy�<�y�<Fy�<ny�<}y�<4y�<�y�<�y�<fy�<=y�<;y�<`   `   xy�<`y�<�y�<�y�<hy�<�y�<ey�<y�<|y�<Uy�<ry�<9y�<Hy�<9y�<ry�<Uy�<|y�<y�<ey�<�y�<hy�<�y�<�y�<`y�<`   `   �y�<{y�<gy�<�y�<Zy�<ly�<uy�<�y�<ny�<ay�<Ky�<y�<�y�<y�<Ky�<ay�<ny�<�y�<uy�<ly�<Zy�<�y�<gy�<{y�<`   `   qy�<Ay�<.y�<�y�<oy�<_y�<^y�<^y�<iy�<�y�<�y�<2y�<�y�<2y�<�y�<�y�<iy�<^y�<^y�<_y�<oy�<�y�<.y�<Ay�<`   `   Iy�<Yy�<dy�<uy�<9y�<]y�<@y�<7y�<zy�<�y�<xy�<+y�<Fy�<+y�<xy�<�y�<zy�<7y�<@y�<]y�<9y�<uy�<dy�<Yy�<`   `   ]y�<�y�<�y�<Oy�<5y�<ay�<ay�<cy�<cy�<<y�<>y�<>y�<py�<>y�<>y�<<y�<cy�<cy�<ay�<ay�<5y�<Oy�<�y�<�y�<`   `   :y�<�y�<my�<�y�<�y�<Jy�<|y�<�y�<Ny�<by�<ty�<qy�<�y�<qy�<ty�<by�<Ny�<�y�<|y�<Jy�<�y�<�y�<my�<�y�<`   `   Sy�<}y�<By�<zy�<ny�<*y�<�y�<}y�<my�<�y�<ry�<Ky�<ay�<Ky�<ry�<�y�<my�<}y�<�y�<*y�<ny�<zy�<By�<}y�<`   `   �y�<�y�<6y�<Sy�<<y�<My�<�y�<Gy�<vy�<7y�<Ay�<Vy�<<y�<Vy�<Ay�<7y�<vy�<Gy�<�y�<My�<<y�<Sy�<6y�<�y�<`   `   Xy�<�y�<Ey�<^y�<Wy�<{y�<�y�<Fy�<�y�<-y�<Vy�<�y�<\y�<�y�<Vy�<-y�<�y�<Fy�<�y�<{y�<Wy�<^y�<Ey�<�y�<`   `   jy�<�y�<Zy�<Gy�<ay�<|y�<vy�<`y�<vy�<*y�<Ey�<~y�<py�<~y�<Ey�<*y�<vy�<`y�<vy�<|y�<ay�<Gy�<Zy�<�y�<`   `   �y�<�y�<cy�<9y�<Wy�<fy�<_y�<Ry�<7y�<5y�<Sy�<{y�<ny�<{y�<Sy�<5y�<7y�<Ry�<_y�<fy�<Wy�<9y�<cy�<�y�<`   `   Dy�<;y�<|y�<_y�<jy�<^y�<cy�<jy�<Gy�<y�<�y�<ny�<2y�<ny�<�y�<y�<Gy�<jy�<cy�<^y�<jy�<_y�<|y�<;y�<`   `   �y�<{y�<�y�<Ty�<�y�<oy�<\y�<ry�<Gy�<py�<]y�<py�<Ry�<py�<]y�<py�<Gy�<ry�<\y�<oy�<�y�<Ty�<�y�<{y�<`   `   yy�<fy�<Yy�<7y�<�y�<ky�<?y�<~y�<Sy�<Ny�<gy�<�y�<y�<�y�<gy�<Ny�<Sy�<~y�<?y�<ky�<�y�<7y�<Yy�<fy�<`   `   -y�<+y�<`y�<`y�<Oy�<:y�<6y�<�y�<xy�<My�<�y�<ky�</y�<ky�<�y�<My�<xy�<�y�<6y�<:y�<Oy�<`y�<`y�<+y�<`   `   �y�<uy�<�y�<py�<y�<^y�<Ly�<ly�<uy�<My�<[y�<,y�<@y�<,y�<[y�<My�<uy�<ly�<Ly�<^y�<y�<py�<�y�<uy�<`   `   �y�<|y�<~y�<^y�<#y�<�y�<Hy�<2y�<iy�<my�<Ly�<Gy�<�y�<Gy�<Ly�<my�<iy�<2y�<Hy�<�y�<#y�<^y�<~y�<|y�<`   `   Ey�<Ty�<vy�<y�<-y�<=y�<Ny�<ay�<Qy�<Dy�<[y�<Xy�<�y�<Xy�<[y�<Dy�<Qy�<ay�<Ny�<=y�<-y�<y�<vy�<Ty�<`   `   xy�<_y�<[y�<�y�<ey�<By�<�y�<�y�<ly�<>y�<ty�<cy�<By�<cy�<ty�<>y�<ly�<�y�<�y�<By�<ey�<�y�<[y�<_y�<`   `   �y�<�y�<z�<�y�<z�<4z�<z�<�y�<�y�<z�<�y�<�y�<z�<�y�<�y�<z�<�y�<�y�<z�<4z�<z�<�y�<z�<�y�<`   `   �y�<z�<	z�<�y�<z�<z�<�y�<�y�< z�<'z�<�y�<�y�<
z�<�y�<�y�<'z�< z�<�y�<�y�<z�<z�<�y�<	z�<z�<`   `   Vz�<z�<�y�<�y�<z�<�y�<�y�<z�<z�<z�<z�<(z�<z�<(z�<z�<z�<z�<z�<�y�<�y�<z�<�y�<�y�<z�<`   `   �y�<�y�<�y�<z�<1z�<%z�<�y�<z�<z�<�y�<�y�<z�<�y�<z�<�y�<�y�<z�<z�<�y�<%z�<1z�<z�<�y�<�y�<`   `   z�<�y�<z�<z�<�y�<�y�<�y�<�y�<�y�<z�<z�<�y�<�y�<�y�<z�<z�<�y�<�y�<�y�<�y�<�y�<z�<z�<�y�<`   `   yz�<z�<�y�<z�<�y�<�y�<�y�<�y�<�y�<�y�<z�<z�<�y�<z�<z�<�y�<�y�<�y�<�y�<�y�<�y�<z�<�y�<z�<`   `   .z�<�y�<�y�<z�<�y�<z�<!z�<�y�<�y�<�y�<�y�<z�<�y�<z�<�y�<�y�<�y�<�y�<!z�<z�<�y�<z�<�y�<�y�<`   `   z�<(z�<z�<�y�<�y�<z�<z�<�y�<z�<�y�<z�<z�<�y�<z�<z�<�y�<z�<�y�<z�<z�<�y�<�y�<z�<(z�<`   `   z�<9z�<+z�<�y�<�y�<z�<z�<z�<z�<,z�<$z�<�y�<z�<�y�<$z�<,z�<z�<z�<z�<z�<�y�<�y�<+z�<9z�<`   `   �y�<�y�<�y�<�y�<z�<z�<z�< z�<�y�<�y�<�y�<�y�<z�<�y�<�y�<�y�<�y�< z�<z�<z�<z�<�y�<�y�<�y�<`   `   .z�<z�<z�<$z�<z�<�y�<�y�<z�<z�<�y�<�y�<z�<z�<z�<�y�<�y�<z�<z�<�y�<�y�<z�<$z�<z�<z�<`   `   z�<�y�<z�<z�<�y�<�y�<�y�<z�<!z�<�y�<z�<#z�<�y�<#z�<z�<�y�<!z�<z�<�y�<�y�<�y�<z�<z�<�y�<`   `   �y�<z�<z�<�y�<�y�<�y�<z�<z�<z�<z�<z�<z�<�y�<z�<z�<z�<z�<z�<z�<�y�<�y�<�y�<z�<z�<`   `   z�<z�<2z�<)z�<%z�<z�<�y�<�y�<z�<z�<�y�<
z�<�y�<
z�<�y�<z�<z�<�y�<�y�<z�<%z�<)z�<2z�<z�<`   `   �y�<�y�<z�<ez�<'z�<�y�<�y�<�y�<z�<z�<�y�<�y�<�y�<�y�<�y�<z�<z�<�y�<�y�<�y�<'z�<ez�<z�<�y�<`   `   z�<�y�<�y�<+z�<�y�<�y�<z�<z�<z�<z�<,z�<z�<�y�<z�<,z�<z�<z�<z�<z�<�y�<�y�<+z�<�y�<�y�<`   `   z�<z�<�y�<z�<z�<"z�<#z�<z�<�y�<�y�<(z�<�y�<�y�<�y�<(z�<�y�<�y�<z�<#z�<"z�<z�<z�<�y�<z�<`   `   �y�<�y�<�y�<z�<�y�<z�<�y�<�y�<�y�<�y�<�y�<�y�<z�<�y�<�y�<�y�<�y�<�y�<�y�<z�<�y�<z�<�y�<�y�<`   `   �y�<�y�<�y�<z�<�y�<z�<�y�<%z�<z�<z�<z�<�y�<Hz�<�y�<z�<z�<z�<%z�<�y�<z�<�y�<z�<�y�<�y�<`   `   
z�< z�<z�<�y�<z�<z�<�y�<Qz�<�y�<z�<6z�<z�<@z�<z�<6z�<z�<�y�<Qz�<�y�<z�<z�<�y�<z�< z�<`   `   Kz�<(z�<z�<�y�<�y�<z�<�y�<#z�<�y�<�y�<�y�<z�<�y�<z�<�y�<�y�<�y�<#z�<�y�<z�<�y�<�y�<z�<(z�<`   `   %z�<�y�<z�<"z�<�y�<z�<+z�<z�<Yz�<z�<�y�<�y�<�y�<�y�<�y�<z�<Yz�<z�<+z�<z�<�y�<"z�<z�<�y�<`   `   z�<�y�<z�<6z�<�y�<
z�<,z�<�y�<Fz�<z�<�y�<z�<�y�<z�<�y�<z�<Fz�<�y�<,z�<
z�<�y�<6z�<z�<�y�<`   `   "z�<�y�<z�<z�<�y�<�y�<z�<�y�<�y�<�y�<�y�<)z�<�y�<)z�<�y�<�y�<�y�<�y�<z�<�y�<�y�<z�<z�<�y�<`   `   z�<�y�<�y�<z�<�y�<�y�<z�<4z�<z�<�y�<z�<�y�<�y�<�y�<z�<�y�<z�<4z�<z�<�y�<�y�<z�<�y�<�y�<`   `   
z�<�y�<�y�<'z�< z�<�y�<�y�<z�<z�<�y�<	z�<z�<�y�<z�<	z�<�y�<z�<z�<�y�<�y�< z�<'z�<�y�<�y�<`   `   z�<(z�<z�<z�<z�<z�<�y�<�y�<z�<�y�<�y�<z�<Vz�<z�<�y�<�y�<z�<�y�<�y�<z�<z�<z�<z�<(z�<`   `   �y�<z�<�y�<�y�<z�<z�<�y�<%z�<1z�<z�<�y�<�y�<�y�<�y�<�y�<z�<1z�<%z�<�y�<z�<z�<�y�<�y�<z�<`   `   �y�<�y�<z�<z�<�y�<�y�<�y�<�y�<�y�<z�<z�<�y�<z�<�y�<z�<z�<�y�<�y�<�y�<�y�<�y�<z�<z�<�y�<`   `   �y�<z�<z�<�y�<�y�<�y�<�y�<�y�<�y�<z�<�y�<z�<yz�<z�<�y�<z�<�y�<�y�<�y�<�y�<�y�<�y�<z�<z�<`   `   �y�<z�<�y�<�y�<�y�<�y�<!z�<z�<�y�<z�<�y�<�y�<.z�<�y�<�y�<z�<�y�<z�<!z�<�y�<�y�<�y�<�y�<z�<`   `   �y�<z�<z�<�y�<z�<�y�<z�<z�<�y�<�y�<z�<(z�<z�<(z�<z�<�y�<�y�<z�<z�<�y�<z�<�y�<z�<z�<`   `   z�<�y�<$z�<,z�<z�<z�<z�<z�<�y�<�y�<+z�<9z�<z�<9z�<+z�<�y�<�y�<z�<z�<z�<z�<,z�<$z�<�y�<`   `   z�<�y�<�y�<�y�<�y�< z�<z�<z�<z�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<z�<z�<z�< z�<�y�<�y�<�y�<�y�<`   `   z�<z�<�y�<�y�<z�<z�<�y�<�y�<z�<$z�<z�<z�<.z�<z�<z�<$z�<z�<�y�<�y�<z�<z�<�y�<�y�<z�<`   `   �y�<#z�<z�<�y�<!z�<z�<�y�<�y�<�y�<z�<z�<�y�<z�<�y�<z�<z�<�y�<�y�<�y�<z�<!z�<�y�<z�<#z�<`   `   �y�<z�<z�<z�<z�<z�<z�<�y�<�y�<�y�<z�<z�<�y�<z�<z�<�y�<�y�<�y�<z�<z�<z�<z�<z�<z�<`   `   �y�<
z�<�y�<z�<z�<�y�<�y�<z�<%z�<)z�<2z�<z�<z�<z�<2z�<)z�<%z�<z�<�y�<�y�<z�<z�<�y�<
z�<`   `   �y�<�y�<�y�<z�<z�<�y�<�y�<�y�<'z�<ez�<z�<�y�<�y�<�y�<z�<ez�<'z�<�y�<�y�<�y�<z�<z�<�y�<�y�<`   `   �y�<z�<,z�<z�<z�<z�<z�<�y�<�y�<+z�<�y�<�y�<z�<�y�<�y�<+z�<�y�<�y�<z�<z�<z�<z�<,z�<z�<`   `   �y�<�y�<(z�<�y�<�y�<z�<#z�<"z�<z�<z�<�y�<z�<z�<z�<�y�<z�<z�<"z�<#z�<z�<�y�<�y�<(z�<�y�<`   `   z�<�y�<�y�<�y�<�y�<�y�<�y�<z�<�y�<z�<�y�<�y�<�y�<�y�<�y�<z�<�y�<z�<�y�<�y�<�y�<�y�<�y�<�y�<`   `   Hz�<�y�<z�<z�<z�<%z�<�y�<z�<�y�<z�<�y�<�y�<�y�<�y�<�y�<z�<�y�<z�<�y�<%z�<z�<z�<z�<�y�<`   `   @z�<z�<6z�<z�<�y�<Qz�<�y�<z�<z�<�y�<z�< z�<
z�< z�<z�<�y�<z�<z�<�y�<Qz�<�y�<z�<6z�<z�<`   `   �y�<z�<�y�<�y�<�y�<#z�<�y�<z�<�y�<�y�<z�<(z�<Kz�<(z�<z�<�y�<�y�<z�<�y�<#z�<�y�<�y�<�y�<z�<`   `   �y�<�y�<�y�<z�<Yz�<z�<+z�<z�<�y�<"z�<z�<�y�<%z�<�y�<z�<"z�<�y�<z�<+z�<z�<Yz�<z�<�y�<�y�<`   `   �y�<z�<�y�<z�<Fz�<�y�<,z�<
z�<�y�<6z�<z�<�y�<z�<�y�<z�<6z�<�y�<
z�<,z�<�y�<Fz�<z�<�y�<z�<`   `   �y�<)z�<�y�<�y�<�y�<�y�<z�<�y�<�y�<z�<z�<�y�<"z�<�y�<z�<z�<�y�<�y�<z�<�y�<�y�<�y�<�y�<)z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   kz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   +z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<
{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<
{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   Tz�<�z�<yz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<yz�<�z�<`   `   �z�<�z�<|z�<�z�<�z�<�z�<�z�<�z�<�z�<xz�<�z�<�z�<�z�<�z�<�z�<xz�<�z�<�z�<�z�<�z�<�z�<�z�<|z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   oz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<|z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<|z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<yz�<�z�<�z�<\z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<){�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<\z�<�z�<�z�<yz�<`   `   �z�<�z�<�z�<lz�<[z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<[z�<lz�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<lz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<lz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   xz�<�z�<�z�<�z�<�z�<�z�<�z�<yz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<yz�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   Ez�<�z�<�z�<�z�<�z�<�z�<�z�<Iz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<Iz�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   {z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<kz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<
{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<+z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<
{�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<yz�<�z�<Tz�<�z�<yz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<xz�<�z�<�z�<�z�<�z�<�z�<�z�<|z�<�z�<�z�<�z�<|z�<�z�<�z�<�z�<�z�<�z�<�z�<xz�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<oz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<|z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<|z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   ){�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<\z�<�z�<�z�<yz�<�z�<yz�<�z�<�z�<\z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<[z�<lz�<�z�<�z�<�z�<�z�<�z�<lz�<[z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<lz�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<lz�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<yz�<�z�<�z�<�z�<�z�<�z�<�z�<xz�<�z�<�z�<�z�<�z�<�z�<�z�<yz�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<Iz�<�z�<�z�<�z�<�z�<�z�<�z�<Ez�<�z�<�z�<�z�<�z�<�z�<�z�<Iz�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �{�<j{�<2{�<{{�<c{�<5{�<?{�<r{�<;{�<a{�<�{�<f{�<V{�<f{�<�{�<a{�<;{�<r{�<?{�<5{�<c{�<{{�<2{�<j{�<`   `   x{�<_{�<>{�<s{�<�{�<p{�<`{�<P{�<T{�<e{�<�{�<|{�<u{�<|{�<�{�<e{�<T{�<P{�<`{�<p{�<�{�<s{�<>{�<_{�<`   `   �z�<H{�<b{�<U{�<y{�<�{�<{{�<V{�<�{�<g{�<?{�<o{�<~{�<o{�<?{�<g{�<�{�<V{�<{{�<�{�<y{�<U{�<b{�<H{�<`   `   b{�<�{�<~{�<]{�<V{�<H{�<O{�<x{�<�{�<j{�<j{�<�{�<}{�<�{�<j{�<j{�<�{�<x{�<O{�<H{�<V{�<]{�<~{�<�{�<`   `   �{�<�{�<v{�<�{�<�{�<M{�<'{�<d{�<j{�<H{�<h{�<i{�<Y{�<i{�<h{�<H{�<j{�<d{�<'{�<M{�<�{�<�{�<v{�<�{�<`   `   A{�<e{�<R{�<P{�<t{�<w{�<[{�<N{�<.{�<7{�<M{�<M{�<�{�<M{�<M{�<7{�<.{�<N{�<[{�<w{�<t{�<P{�<R{�<e{�<`   `   w{�<�{�<e{�<={�<?{�<^{�<�{�<b{�<.{�<�{�<�{�<k{�<�{�<k{�<�{�<�{�<.{�<b{�<�{�<^{�<?{�<={�<e{�<�{�<`   `   �{�<�{�<W{�<�{�<j{�<[{�<�{�<n{�<G{�<�{�<u{�< {�<f{�< {�<u{�<�{�<G{�<n{�<�{�<[{�<j{�<�{�<W{�<�{�<`   `   �{�<G{�<B{�<�{�<I{�<X{�<n{�<c{�<q{�<W{�<d{�<<{�<L{�<<{�<d{�<W{�<q{�<c{�<n{�<X{�<I{�<�{�<B{�<G{�<`   `   �{�<p{�<j{�<�{�<8{�<j{�<c{�<[{�<�{�<Y{�<�{�<�{�<M{�<�{�<�{�<Y{�<�{�<[{�<c{�<j{�<8{�<�{�<j{�<p{�<`   `   ~{�<�{�<`{�<b{�<o{�<�{�<�{�<s{�<y{�<O{�<m{�<X{�<1{�<X{�<m{�<O{�<y{�<s{�<�{�<�{�<o{�<b{�<`{�<�{�<`   `   n{�<�{�<Z{�<\{�<R{�<P{�<g{�<o{�<�{�<�{�<^{�<^{�<�{�<^{�<^{�<�{�<�{�<o{�<g{�<P{�<R{�<\{�<Z{�<�{�<`   `   W{�<\{�<g{�<�{�<a{�<N{�<H{�<g{�<x{�<�{�<p{�<;{�<x{�<;{�<p{�<�{�<x{�<g{�<H{�<N{�<a{�<�{�<g{�<\{�<`   `   o{�<a{�<e{�<�{�<�{�<|{�<@{�<�{�<]{�<F{�<s{�<{�<.{�<{�<s{�<F{�<]{�<�{�<@{�<|{�<�{�<�{�<e{�<a{�<`   `   q{�<�{�<�{�<|{�<�{�<u{�<?{�<�{�<s{�<p{�<�{�<^{�<h{�<^{�<�{�<p{�<s{�<�{�<?{�<u{�<�{�<|{�<�{�<�{�<`   `   -{�<Z{�<�{�<{�<�{�<`{�<a{�<i{�<T{�<�{�<�{�<q{�<S{�<q{�<�{�<�{�<T{�<i{�<a{�<`{�<�{�<{�<�{�<Z{�<`   `   4{�<={�<p{�<q{�<l{�<;{�<i{�<X{�<K{�<^{�<a{�<v{�<{�<v{�<a{�<^{�<K{�<X{�<i{�<;{�<l{�<q{�<p{�<={�<`   `   A{�<N{�<�{�<d{�<�{�<c{�<i{�<�{�<�{�<d{�<`{�<�{�<{�<�{�<`{�<d{�<�{�<�{�<i{�<c{�<�{�<d{�<�{�<N{�<`   `   R{�<j{�<�{�<G{�<�{�<�{�<M{�<M{�<~{�<W{�<`{�<�{�<G{�<�{�<`{�<W{�<~{�<M{�<M{�<�{�<�{�<G{�<�{�<j{�<`   `   m{�<s{�<_{�<[{�<v{�<|{�<d{�<P{�<�{�<\{�<W{�<�{�<a{�<�{�<W{�<\{�<�{�<P{�<d{�<|{�<v{�<[{�<_{�<s{�<`   `   m{�<�{�<_{�<�{�<�{�<n{�<�{�<�{�<�{�<�{�<w{�<j{�<d{�<j{�<w{�<�{�<�{�<�{�<�{�<n{�<�{�<�{�<_{�<�{�<`   `   �{�<�{�<T{�<g{�<a{�<:{�<z{�<�{�<O{�<e{�<�{�<Z{�<p{�<Z{�<�{�<e{�<O{�<�{�<z{�<:{�<a{�<g{�<T{�<�{�<`   `   }{�<o{�<G{�<j{�<|{�<S{�<h{�<�{�<R{�<f{�<s{�<{�<I{�<{�<s{�<f{�<R{�<�{�<h{�<S{�<|{�<j{�<G{�<o{�<`   `   L{�<?{�<t{�<�{�<}{�<�{�<^{�<�{�<y{�<�{�<R{�<${�<�{�<${�<R{�<�{�<y{�<�{�<^{�<�{�<}{�<�{�<t{�<?{�<`   `   V{�<f{�<�{�<a{�<;{�<r{�<?{�<5{�<c{�<{{�<2{�<j{�<�{�<j{�<2{�<{{�<c{�<5{�<?{�<r{�<;{�<a{�<�{�<f{�<`   `   u{�<|{�<�{�<e{�<T{�<P{�<`{�<p{�<�{�<s{�<>{�<_{�<x{�<_{�<>{�<s{�<�{�<p{�<`{�<P{�<T{�<e{�<�{�<|{�<`   `   ~{�<o{�<?{�<g{�<�{�<V{�<{{�<�{�<y{�<U{�<b{�<H{�<�z�<H{�<b{�<U{�<y{�<�{�<{{�<V{�<�{�<g{�<?{�<o{�<`   `   }{�<�{�<j{�<j{�<�{�<x{�<O{�<H{�<V{�<]{�<~{�<�{�<b{�<�{�<~{�<]{�<V{�<H{�<O{�<x{�<�{�<j{�<j{�<�{�<`   `   Y{�<i{�<h{�<H{�<j{�<d{�<'{�<M{�<�{�<�{�<v{�<�{�<�{�<�{�<v{�<�{�<�{�<M{�<'{�<d{�<j{�<H{�<h{�<i{�<`   `   �{�<M{�<M{�<7{�<.{�<N{�<[{�<w{�<t{�<P{�<R{�<e{�<A{�<e{�<R{�<P{�<t{�<w{�<[{�<N{�<.{�<7{�<M{�<M{�<`   `   �{�<k{�<�{�<�{�<.{�<b{�<�{�<^{�<?{�<={�<e{�<�{�<w{�<�{�<e{�<={�<?{�<^{�<�{�<b{�<.{�<�{�<�{�<k{�<`   `   f{�< {�<u{�<�{�<G{�<n{�<�{�<[{�<j{�<�{�<W{�<�{�<�{�<�{�<W{�<�{�<j{�<[{�<�{�<n{�<G{�<�{�<u{�< {�<`   `   L{�<<{�<d{�<W{�<q{�<c{�<n{�<X{�<I{�<�{�<B{�<G{�<�{�<G{�<B{�<�{�<I{�<X{�<n{�<c{�<q{�<W{�<d{�<<{�<`   `   M{�<�{�<�{�<Y{�<�{�<[{�<c{�<j{�<8{�<�{�<j{�<p{�<�{�<p{�<j{�<�{�<8{�<j{�<c{�<[{�<�{�<Y{�<�{�<�{�<`   `   1{�<X{�<m{�<O{�<y{�<s{�<�{�<�{�<o{�<b{�<`{�<�{�<~{�<�{�<`{�<b{�<o{�<�{�<�{�<s{�<y{�<O{�<m{�<X{�<`   `   �{�<^{�<^{�<�{�<�{�<o{�<g{�<P{�<R{�<\{�<Z{�<�{�<n{�<�{�<Z{�<\{�<R{�<P{�<g{�<o{�<�{�<�{�<^{�<^{�<`   `   x{�<;{�<p{�<�{�<x{�<g{�<H{�<N{�<a{�<�{�<g{�<\{�<W{�<\{�<g{�<�{�<a{�<N{�<H{�<g{�<x{�<�{�<p{�<;{�<`   `   .{�<{�<s{�<F{�<]{�<�{�<@{�<|{�<�{�<�{�<e{�<a{�<o{�<a{�<e{�<�{�<�{�<|{�<@{�<�{�<]{�<F{�<s{�<{�<`   `   h{�<^{�<�{�<p{�<s{�<�{�<?{�<u{�<�{�<|{�<�{�<�{�<q{�<�{�<�{�<|{�<�{�<u{�<?{�<�{�<s{�<p{�<�{�<^{�<`   `   S{�<q{�<�{�<�{�<T{�<i{�<a{�<`{�<�{�<{�<�{�<Z{�<-{�<Z{�<�{�<{�<�{�<`{�<a{�<i{�<T{�<�{�<�{�<q{�<`   `   {�<v{�<a{�<^{�<K{�<X{�<i{�<;{�<l{�<q{�<p{�<={�<4{�<={�<p{�<q{�<l{�<;{�<i{�<X{�<K{�<^{�<a{�<v{�<`   `   {�<�{�<`{�<d{�<�{�<�{�<i{�<c{�<�{�<d{�<�{�<N{�<A{�<N{�<�{�<d{�<�{�<c{�<i{�<�{�<�{�<d{�<`{�<�{�<`   `   G{�<�{�<`{�<W{�<~{�<M{�<M{�<�{�<�{�<G{�<�{�<j{�<R{�<j{�<�{�<G{�<�{�<�{�<M{�<M{�<~{�<W{�<`{�<�{�<`   `   a{�<�{�<W{�<\{�<�{�<P{�<d{�<|{�<v{�<[{�<_{�<s{�<m{�<s{�<_{�<[{�<v{�<|{�<d{�<P{�<�{�<\{�<W{�<�{�<`   `   d{�<j{�<w{�<�{�<�{�<�{�<�{�<n{�<�{�<�{�<_{�<�{�<m{�<�{�<_{�<�{�<�{�<n{�<�{�<�{�<�{�<�{�<w{�<j{�<`   `   p{�<Z{�<�{�<e{�<O{�<�{�<z{�<:{�<a{�<g{�<T{�<�{�<�{�<�{�<T{�<g{�<a{�<:{�<z{�<�{�<O{�<e{�<�{�<Z{�<`   `   I{�<{�<s{�<f{�<R{�<�{�<h{�<S{�<|{�<j{�<G{�<o{�<}{�<o{�<G{�<j{�<|{�<S{�<h{�<�{�<R{�<f{�<s{�<{�<`   `   �{�<${�<R{�<�{�<y{�<�{�<^{�<�{�<}{�<�{�<t{�<?{�<L{�<?{�<t{�<�{�<}{�<�{�<^{�<�{�<y{�<�{�<R{�<${�<`   `   �{�<3|�<G|�<�{�<6|�<\|�<N|�<#|�<|�<6|�<|�<"|�<�|�<"|�<|�<6|�<|�<#|�<N|�<\|�<6|�<�{�<G|�<3|�<`   `   |�<h|�<f|�<3|�<|�<0|�<'|�<*|�<i|�<E|�< |�<|�<|�<|�< |�<E|�<i|�<*|�<'|�<0|�<|�<3|�<f|�<h|�<`   `   p|�<c|�<E|�<7|�<|�<)|�<4|�<0|�<<|�<1|�<C|�<,|�<|�<,|�<C|�<1|�<<|�<0|�<4|�<)|�<|�<7|�<E|�<c|�<`   `   A|�<|�< |�<|�<9|�<`|�<H|�<,|�<|�<|�<=|�<4|�<5|�<4|�<=|�<|�<|�<,|�<H|�<`|�<9|�<|�< |�<|�<`   `   D|�<|�<>|�<C|�<!|�<M|�<*|�<H|�<B|�<H|�<[|�<(|�<|�<(|�<[|�<H|�<B|�<H|�<*|�<M|�<!|�<C|�<>|�<|�<`   `   `|�<|�<K|�<O|�<|�<F|�<4|�<l|�<^|�<C|�<a|�<)|�<�{�<)|�<a|�<C|�<^|�<l|�<4|�<F|�<|�<O|�<K|�<|�<`   `   X|�<�{�<!|�<?|�<&|�<?|�<|�<N|�<+|�<|�<%|�<.|�<?|�<.|�<%|�<|�<+|�<N|�<|�<?|�<&|�<?|�<!|�<�{�<`   `   |�<	|�<P|�<A|�<9|�<C|�<
|�<7|�<B|�<;|�<|�<,|�<[|�<,|�<|�<;|�<B|�<7|�<
|�<C|�<9|�<A|�<P|�<	|�<`   `   |�<5|�<h|�<|�<|�<`|�<-|�<4|�<W|�<R|�<8|�<T|�<S|�<T|�<8|�<R|�<W|�<4|�<-|�<`|�<|�<|�<h|�<5|�<`   `   &|�<$|�<)|�<|�<:|�<O|�<.|�<+|�<,|�<|�<|�<e|�<?|�<e|�<|�<|�<,|�<+|�<.|�<O|�<:|�<|�<)|�<$|�<`   `   |�<|�<&|�<c|�<v|�<|�<|�<3|�<8|�<|�<|�<7|�<�{�<7|�<|�<|�<8|�<3|�<|�<|�<v|�<c|�<&|�<|�<`   `   |�<@|�<;|�<S|�<*|�<|�<7|�<|�<7|�<-|�<7|�<W|�<&|�<W|�<7|�<-|�<7|�<|�<7|�<|�<*|�<S|�<;|�<@|�<`   `   |�<F|�<|�<|�<�{�<]|�<�|�<|�</|�<#|�<K|�<f|�<?|�<f|�<K|�<#|�</|�<|�<�|�<]|�<�{�<|�<|�<F|�<`   `   |�<b|�<%|�<|�<|�<A|�<M|�<|�<@|�< |�<@|�<D|�<+|�<D|�<@|�< |�<@|�<|�<M|�<A|�<|�<|�<%|�<b|�<`   `   |�<=|�<|�<|�<|�<�{�<|�<|�<B|�<|�<|�<D|�<\|�<D|�<|�<|�<B|�<|�<|�<�{�<|�<|�<|�<=|�<`   `   S|�<|�<|�<|�<|�<<|�<n|�<E|�<J|�<3|�<|�<8|�<S|�<8|�<|�<3|�<J|�<E|�<n|�<<|�<|�<|�<|�<|�<`   `   �|�<N|�<8|�<:|�<|�<K|�<m|�<|�<|�<O|�<$|�<?|�</|�<?|�<$|�<O|�<|�<|�<m|�<K|�<|�<:|�<8|�<N|�<`   `   �|�<|�<3|�<1|�<B|�<2|�<+|�<"|�<
|�<<|�<|�<C|�<C|�<C|�<|�<<|�<
|�<"|�<+|�<2|�<B|�<1|�<3|�<|�<`   `   $|�<|�<A|�<|�<5|�< |�< |�<g|�<J|�<B|�<|�<3|�<C|�<3|�<|�<B|�<J|�<g|�< |�< |�<5|�<|�<A|�<|�<`   `   :|�<=|�<J|�<|�<|�<%|�<|�<1|�<|�<-|�<P|�<0|�<#|�<0|�<P|�<-|�<|�<1|�<|�<%|�<|�<|�<J|�<=|�<`   `    |�<|�<|�<A|�<|�<<|�<%|�<|�<�{�<|�<>|�<|�<4|�<|�<>|�<|�<�{�<|�<%|�<<|�<|�<A|�<|�<|�<`   `   |�<|�<5|�<N|�<|�<:|�<
|�<2|�<T|�<%|�<|�<|�<}|�<|�<|�<%|�<T|�<2|�<
|�<:|�<|�<N|�<5|�<|�<`   `   #|�<|�<H|�<W|�<|�<a|�<|�<�{�<A|�<8|�<H|�<P|�<�|�<P|�<H|�<8|�<A|�<�{�<|�<a|�<|�<W|�<H|�<|�<`   `   {|�<|�<&|�<H|�<�{�<U|�<E|�<|�<|�<
|�<l|�<j|�<'|�<j|�<l|�<
|�<|�<|�<E|�<U|�<�{�<H|�<&|�<|�<`   `   �|�<"|�<|�<6|�<|�<#|�<N|�<\|�<6|�<�{�<G|�<3|�<�{�<3|�<G|�<�{�<6|�<\|�<N|�<#|�<|�<6|�<|�<"|�<`   `   |�<|�< |�<E|�<i|�<*|�<'|�<0|�<|�<3|�<f|�<h|�<|�<h|�<f|�<3|�<|�<0|�<'|�<*|�<i|�<E|�< |�<|�<`   `   |�<,|�<C|�<1|�<<|�<0|�<4|�<)|�<|�<7|�<E|�<c|�<p|�<c|�<E|�<7|�<|�<)|�<4|�<0|�<<|�<1|�<C|�<,|�<`   `   5|�<4|�<=|�<|�<|�<,|�<H|�<`|�<9|�<|�< |�<|�<A|�<|�< |�<|�<9|�<`|�<H|�<,|�<|�<|�<=|�<4|�<`   `   |�<(|�<[|�<H|�<B|�<H|�<*|�<M|�<!|�<C|�<>|�<|�<D|�<|�<>|�<C|�<!|�<M|�<*|�<H|�<B|�<H|�<[|�<(|�<`   `   �{�<)|�<a|�<C|�<^|�<l|�<4|�<F|�<|�<O|�<K|�<|�<`|�<|�<K|�<O|�<|�<F|�<4|�<l|�<^|�<C|�<a|�<)|�<`   `   ?|�<.|�<%|�<|�<+|�<N|�<|�<?|�<&|�<?|�<!|�<�{�<X|�<�{�<!|�<?|�<&|�<?|�<|�<N|�<+|�<|�<%|�<.|�<`   `   [|�<,|�<|�<;|�<B|�<7|�<
|�<C|�<9|�<A|�<P|�<	|�<|�<	|�<P|�<A|�<9|�<C|�<
|�<7|�<B|�<;|�<|�<,|�<`   `   S|�<T|�<8|�<R|�<W|�<4|�<-|�<`|�<|�<|�<h|�<5|�<|�<5|�<h|�<|�<|�<`|�<-|�<4|�<W|�<R|�<8|�<T|�<`   `   ?|�<e|�<|�<|�<,|�<+|�<.|�<O|�<:|�<|�<)|�<$|�<&|�<$|�<)|�<|�<:|�<O|�<.|�<+|�<,|�<|�<|�<e|�<`   `   �{�<7|�<|�<|�<8|�<3|�<|�<|�<v|�<c|�<&|�<|�<|�<|�<&|�<c|�<v|�<|�<|�<3|�<8|�<|�<|�<7|�<`   `   &|�<W|�<7|�<-|�<7|�<|�<7|�<|�<*|�<S|�<;|�<@|�<|�<@|�<;|�<S|�<*|�<|�<7|�<|�<7|�<-|�<7|�<W|�<`   `   ?|�<f|�<K|�<#|�</|�<|�<�|�<]|�<�{�<|�<|�<F|�<|�<F|�<|�<|�<�{�<]|�<�|�<|�</|�<#|�<K|�<f|�<`   `   +|�<D|�<@|�< |�<@|�<|�<M|�<A|�<|�<|�<%|�<b|�<|�<b|�<%|�<|�<|�<A|�<M|�<|�<@|�< |�<@|�<D|�<`   `   \|�<D|�<|�<|�<B|�<|�<|�<�{�<|�<|�<|�<=|�<|�<=|�<|�<|�<|�<�{�<|�<|�<B|�<|�<|�<D|�<`   `   S|�<8|�<|�<3|�<J|�<E|�<n|�<<|�<|�<|�<|�<|�<S|�<|�<|�<|�<|�<<|�<n|�<E|�<J|�<3|�<|�<8|�<`   `   /|�<?|�<$|�<O|�<|�<|�<m|�<K|�<|�<:|�<8|�<N|�<�|�<N|�<8|�<:|�<|�<K|�<m|�<|�<|�<O|�<$|�<?|�<`   `   C|�<C|�<|�<<|�<
|�<"|�<+|�<2|�<B|�<1|�<3|�<|�<�|�<|�<3|�<1|�<B|�<2|�<+|�<"|�<
|�<<|�<|�<C|�<`   `   C|�<3|�<|�<B|�<J|�<g|�< |�< |�<5|�<|�<A|�<|�<$|�<|�<A|�<|�<5|�< |�< |�<g|�<J|�<B|�<|�<3|�<`   `   #|�<0|�<P|�<-|�<|�<1|�<|�<%|�<|�<|�<J|�<=|�<:|�<=|�<J|�<|�<|�<%|�<|�<1|�<|�<-|�<P|�<0|�<`   `   4|�<|�<>|�<|�<�{�<|�<%|�<<|�<|�<A|�<|�<|�< |�<|�<|�<A|�<|�<<|�<%|�<|�<�{�<|�<>|�<|�<`   `   }|�<|�<|�<%|�<T|�<2|�<
|�<:|�<|�<N|�<5|�<|�<|�<|�<5|�<N|�<|�<:|�<
|�<2|�<T|�<%|�<|�<|�<`   `   �|�<P|�<H|�<8|�<A|�<�{�<|�<a|�<|�<W|�<H|�<|�<#|�<|�<H|�<W|�<|�<a|�<|�<�{�<A|�<8|�<H|�<P|�<`   `   '|�<j|�<l|�<
|�<|�<|�<E|�<U|�<�{�<H|�<&|�<|�<{|�<|�<&|�<H|�<�{�<U|�<E|�<|�<|�<
|�<l|�<j|�<`   `   �|�<}�<�|�< }�<;}�<!}�<}�<�|�<<}�<
}�<}�<}�<�|�<}�<}�<
}�<<}�<�|�<}�<!}�<;}�< }�<�|�<}�<`   `   }�<�|�<�|�<}�<�|�<�|�<}�<}�<}�<�|�<}�<}�<�|�<}�<}�<�|�<}�<}�<}�<�|�<�|�<}�<�|�<�|�<`   `   }�<�|�<�|�<3}�<}�<�|�<�|�<}�<�|�<�|�<8}�< }�<}�< }�<8}�<�|�<�|�<}�<�|�<�|�<}�<3}�<�|�<�|�<`   `   �|�<
}�<}�<}�<+}�<�|�<	}�<}�<�|�<&}�<�|�<�|�<"}�<�|�<�|�<&}�<�|�<}�<	}�<�|�<+}�<}�<}�<
}�<`   `   �|�<#}�<&}�<�|�<�|�<�|�<}�<�|�<�|�<	}�<�|�<}�<j}�<}�<�|�<	}�<�|�<�|�<}�<�|�<�|�<�|�<&}�<#}�<`   `   }�<}�<"}�<�|�<}�<}�<�|�<�|�<}�<}�<�|�<6}�<!}�<6}�<�|�<}�<}�<�|�<�|�<}�<}�<�|�<"}�<}�<`   `   )}�< }�<}�<}�<2}�<}�<�|�<�|�<}�< }�<�|�<}�<�|�<}�<�|�< }�<}�<�|�<�|�<}�<2}�<}�<}�< }�<`   `    }�<�|�<}�<�|�<}�<�|�<�|�<}�<�|�<�|�<}�<5}�<�|�<5}�<}�<�|�<�|�<}�<�|�<�|�<}�<�|�<}�<�|�<`   `   }�<}�<}�<�|�</}�<�|�<}�<}�<�|�<}�<�|�<�|�<�|�<�|�<�|�<}�<�|�<}�<}�<�|�</}�<�|�<}�<}�<`   `   .}�<}�<}�<�|�<}�<�|�<}�<}�<�|�<E}�<�|�<�|�<�|�<�|�<�|�<E}�<�|�<}�<}�<�|�<}�<�|�<}�<}�<`   `   !}�<�|�<}�<�|�<�|�<�|�<(}�<%}�<}�<y}�<&}�<}�<9}�<}�<&}�<y}�<}�<%}�<(}�<�|�<�|�<�|�<}�<�|�<`   `   .}�<}�<}�<�|�<}�< }�<}�<}�<�|�<}�<}�<�|�<�|�<�|�<}�<}�<�|�<}�<}�< }�<}�<�|�<}�<}�<`   `   }�< }�<�|�<'}�<3}�<}�<�|�<�|�<}�<�|�<�|�<�|�<�|�<�|�<�|�<�|�<}�<�|�<�|�<}�<3}�<'}�<�|�< }�<`   `   �|�<}�<�|�<.}�<}�<�|�<}�<
}�<<}�<,}�<}�<}�<}�<}�<}�<,}�<<}�<
}�<}�<�|�<}�<.}�<�|�<}�<`   `   �|�<%}�<
}�<%}�<}�<}�<9}�<�|�<�|�<
}�<}�<�|�<�|�<�|�<}�<
}�<�|�<�|�<9}�<}�<}�<%}�<
}�<%}�<`   `   �|�<�|�< }�<"}�<'}�<%}�<�|�<�|�<}�<�|�<�|�<�|�<�|�<�|�<�|�<�|�<}�<�|�<�|�<%}�<'}�<"}�< }�<�|�<`   `   �|�<�|�<5}�<}�<}�<�|�<�|�<}�<>}�<"}�<}�<}�<}�<}�<}�<"}�<>}�<}�<�|�<�|�<}�<}�<5}�<�|�<`   `   �|�<�|�<}�<�|�<}�<�|�<�|�<}�<�|�<}�<}�<�|�<}�<�|�<}�<}�<�|�<}�<�|�<�|�<}�<�|�<}�<�|�<`   `   }�<}�<}�<}�< }�<�|�<*}�< }�<�|�<#}�<�|�<�|�<}�<�|�<�|�<#}�<�|�< }�<*}�<�|�< }�<}�<}�<}�<`   `   }�<}�<}�<-}�<}�<}�<}�<}�<}�<&}�<}�<�|�<}�<�|�<}�<&}�<}�<}�<}�<}�<}�<-}�<}�<}�<`   `   }�<}�<�|�<�|�<}�<"}�<�|�<�|�<	}�<}�</}�<}�<"}�<}�</}�<}�<	}�<�|�<�|�<"}�<}�<�|�<�|�<}�<`   `   }�<0}�<}�<�|�<}�<,}�<}�<}�<'}�<}�<&}�<�|�<�|�<�|�<&}�<}�<'}�<}�<}�<,}�<}�<�|�<}�<0}�<`   `   �|�<$}�<}�<�|�<}�<}�<}�<}�<}�<�|�<�|�<�|�<�|�<�|�<�|�<�|�<}�<}�<}�<}�<}�<�|�<}�<$}�<`   `   �|�<%}�<}�<�|�<}�<�|�<�|�<�|�<}�<�|�<�|�<}�<�|�<}�<�|�<�|�<}�<�|�<�|�<�|�<}�<�|�<}�<%}�<`   `   �|�<}�<}�<
}�<<}�<�|�<}�<!}�<;}�< }�<�|�<}�<�|�<}�<�|�< }�<;}�<!}�<}�<�|�<<}�<
}�<}�<}�<`   `   �|�<}�<}�<�|�<}�<}�<}�<�|�<�|�<}�<�|�<�|�<}�<�|�<�|�<}�<�|�<�|�<}�<}�<}�<�|�<}�<}�<`   `   }�< }�<8}�<�|�<�|�<}�<�|�<�|�<}�<3}�<�|�<�|�<}�<�|�<�|�<3}�<}�<�|�<�|�<}�<�|�<�|�<8}�< }�<`   `   "}�<�|�<�|�<&}�<�|�<}�<	}�<�|�<+}�<}�<}�<
}�<�|�<
}�<}�<}�<+}�<�|�<	}�<}�<�|�<&}�<�|�<�|�<`   `   j}�<}�<�|�<	}�<�|�<�|�<}�<�|�<�|�<�|�<&}�<#}�<�|�<#}�<&}�<�|�<�|�<�|�<}�<�|�<�|�<	}�<�|�<}�<`   `   !}�<6}�<�|�<}�<}�<�|�<�|�<}�<}�<�|�<"}�<}�<}�<}�<"}�<�|�<}�<}�<�|�<�|�<}�<}�<�|�<6}�<`   `   �|�<}�<�|�< }�<}�<�|�<�|�<}�<2}�<}�<}�< }�<)}�< }�<}�<}�<2}�<}�<�|�<�|�<}�< }�<�|�<}�<`   `   �|�<5}�<}�<�|�<�|�<}�<�|�<�|�<}�<�|�<}�<�|�< }�<�|�<}�<�|�<}�<�|�<�|�<}�<�|�<�|�<}�<5}�<`   `   �|�<�|�<�|�<}�<�|�<}�<}�<�|�</}�<�|�<}�<}�<}�<}�<}�<�|�</}�<�|�<}�<}�<�|�<}�<�|�<�|�<`   `   �|�<�|�<�|�<E}�<�|�<}�<}�<�|�<}�<�|�<}�<}�<.}�<}�<}�<�|�<}�<�|�<}�<}�<�|�<E}�<�|�<�|�<`   `   9}�<}�<&}�<y}�<}�<%}�<(}�<�|�<�|�<�|�<}�<�|�<!}�<�|�<}�<�|�<�|�<�|�<(}�<%}�<}�<y}�<&}�<}�<`   `   �|�<�|�<}�<}�<�|�<}�<}�< }�<}�<�|�<}�<}�<.}�<}�<}�<�|�<}�< }�<}�<}�<�|�<}�<}�<�|�<`   `   �|�<�|�<�|�<�|�<}�<�|�<�|�<}�<3}�<'}�<�|�< }�<}�< }�<�|�<'}�<3}�<}�<�|�<�|�<}�<�|�<�|�<�|�<`   `   }�<}�<}�<,}�<<}�<
}�<}�<�|�<}�<.}�<�|�<}�<�|�<}�<�|�<.}�<}�<�|�<}�<
}�<<}�<,}�<}�<}�<`   `   �|�<�|�<}�<
}�<�|�<�|�<9}�<}�<}�<%}�<
}�<%}�<�|�<%}�<
}�<%}�<}�<}�<9}�<�|�<�|�<
}�<}�<�|�<`   `   �|�<�|�<�|�<�|�<}�<�|�<�|�<%}�<'}�<"}�< }�<�|�<�|�<�|�< }�<"}�<'}�<%}�<�|�<�|�<}�<�|�<�|�<�|�<`   `   }�<}�<}�<"}�<>}�<}�<�|�<�|�<}�<}�<5}�<�|�<�|�<�|�<5}�<}�<}�<�|�<�|�<}�<>}�<"}�<}�<}�<`   `   }�<�|�<}�<}�<�|�<}�<�|�<�|�<}�<�|�<}�<�|�<�|�<�|�<}�<�|�<}�<�|�<�|�<}�<�|�<}�<}�<�|�<`   `   }�<�|�<�|�<#}�<�|�< }�<*}�<�|�< }�<}�<}�<}�<}�<}�<}�<}�< }�<�|�<*}�< }�<�|�<#}�<�|�<�|�<`   `   }�<�|�<}�<&}�<}�<}�<}�<}�<}�<-}�<}�<}�<}�<}�<}�<-}�<}�<}�<}�<}�<}�<&}�<}�<�|�<`   `   "}�<}�</}�<}�<	}�<�|�<�|�<"}�<}�<�|�<�|�<}�<}�<}�<�|�<�|�<}�<"}�<�|�<�|�<	}�<}�</}�<}�<`   `   �|�<�|�<&}�<}�<'}�<}�<}�<,}�<}�<�|�<}�<0}�<}�<0}�<}�<�|�<}�<,}�<}�<}�<'}�<}�<&}�<�|�<`   `   �|�<�|�<�|�<�|�<}�<}�<}�<}�<}�<�|�<}�<$}�<�|�<$}�<}�<�|�<}�<}�<}�<}�<}�<�|�<�|�<�|�<`   `   �|�<}�<�|�<�|�<}�<�|�<�|�<�|�<}�<�|�<}�<%}�<�|�<%}�<}�<�|�<}�<�|�<�|�<�|�<}�<�|�<�|�<}�<`   `   G~�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<`   `   ~�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<-~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<-~�<�}�<�}�<�}�<�}�<`   `   �}�<~�<~�<�}�<~�<�}�<�}�<~�<)~�<%~�<�}�<�}�<�}�<�}�<�}�<%~�<)~�<~�<�}�<�}�<~�<�}�<~�<~�<`   `   �}�<�}�<�}�<�}�<"~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<"~�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<`   `   �}�<~�<�}�<�}�<�}�<�}�<"~�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<"~�<�}�<�}�<�}�<�}�<~�<`   `   �}�<~�<�}�<�}�<�}�<�}�<-~�<�}�<�}�<�}�<�}�<~�<
~�<~�<�}�<�}�<�}�<�}�<-~�<�}�<�}�<�}�<�}�<~�<`   `   �}�<�}�<�}�<~�<~�<�}�<~�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<~�<�}�<~�<~�<�}�<�}�<`   `   �}�<�}�<�}�<~�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<~�<�}�<�}�<`   `   �}�<�}�<~�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<~�<�}�<`   `   �}�<�}�<~�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<~�<�}�<`   `   ~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<~�<~�<~�<~�<~�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<~�<�}�<�}�<�}�<~�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<`   `   ~�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<!~�<~�<~�<~�<!~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<`   `   �}�<	~�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<	~�<`   `   ~�<-~�<�}�<�}�<�}�<~�<~�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<~�<~�<�}�<�}�<�}�<-~�<`   `   �}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<~�<�}�<~�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<`   `   �}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�< ~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�< ~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<
~�<~�<�}�<~�<
~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<~�<�}�<~�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<~�<�}�<~�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<
~�<�}�<~�<�}�<�}�<~�<�}�<�}�<~�<�}�<�}�<~�<�}�<�}�<~�<�}�<
~�<�}�<�}�<�}�<`   `   �}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<G~�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   ~�<�}�<�}�<�}�<�}�<�}�<�}�<-~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<-~�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<%~�<)~�<~�<�}�<�}�<~�<�}�<~�<~�<�}�<~�<~�<�}�<~�<�}�<�}�<~�<)~�<%~�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<"~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<"~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<~�<�}�<�}�<"~�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<"~�<�}�<�}�<~�<�}�<�}�<`   `   
~�<~�<�}�<�}�<�}�<�}�<-~�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<-~�<�}�<�}�<�}�<�}�<~�<`   `   �}�<~�<�}�<�}�<�}�<�}�<~�<�}�<~�<~�<�}�<�}�<�}�<�}�<�}�<~�<~�<�}�<~�<�}�<�}�<�}�<�}�<~�<`   `   �}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<~�<�}�<�}�<�}�<�}�<�}�<~�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<`   `   ~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<~�<�}�<�}�<�}�<~�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<~�<�}�<�}�<�}�<~�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<`   `   ~�<~�<~�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<~�<~�<`   `   ~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<~�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<~�<�}�<`   `   ~�<~�<!~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<~�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<!~�<~�<`   `   �}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<	~�<�}�<	~�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<�}�<~�<~�<~�<�}�<�}�<�}�<-~�<~�<-~�<�}�<�}�<�}�<~�<~�<~�<�}�<�}�<�}�<�}�<`   `   �}�<~�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<~�<`   `   �}�<�}�<�}�<�}�< ~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�< ~�<�}�<�}�<�}�<`   `   �}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<`   `   �}�<~�<
~�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<
~�<~�<`   `   �}�<�}�<�}�<�}�<�}�<~�<~�<�}�<~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<~�<�}�<~�<~�<�}�<�}�<�}�<�}�<`   `   ~�<�}�<�}�<~�<�}�<�}�<~�<�}�<
~�<�}�<�}�<�}�<�}�<�}�<�}�<�}�<
~�<�}�<~�<�}�<�}�<~�<�}�<�}�<`   `   Y~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<|~�<�~�<�<�~�<�<�~�<|~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �<�~�<�~�<	�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<	�<�~�<�~�<`   `   �<�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<5�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�<�~�<	�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<	�<�~�<�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<	�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�<�~�<�~�<�~�<�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<	�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �<�~�<�~�<�~�<�~�<�<"�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<"�<�<�~�<�~�<�~�<�~�<`   `   �~�<�~�< �<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�< �<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<`   `   �~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<`   `   �~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�<�<�~�<�~�<�~�<�~�<�~�<�<�<�~�<�~�<�~�<�~�<�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<
�<�~�<�~�<�~�<�~�<�~�<
�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<Y~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<`   `   �<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�<�~�<|~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<|~�<�~�<�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<	�<�~�<�~�<�<�~�<�~�<	�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�<�<�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<`   `   5�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<	�<�~�<�<�~�<�~�<�~�<�~�<�~�<�<�~�<	�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<	�<�~�<	�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<"�<�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�<"�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�< �<�~�<�~�<�~�< �<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�<�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�<�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<`   `   �~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<`   `   �~�<�~�<�~�<
�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<
�<�~�<�~�<`   `   �~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   �~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<`   `   Z��<
��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<
��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��< ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��< ��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<%��<��<��<��<%��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<2��<��<��<-��<��<��<��<-��<��<��<2��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<.��<��<��<��<��<��<��<��<��<��<��<��<`   `   Y�<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��</��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `    ��<��<��<��<��<��<��<��<��<��<��<!��<��<!��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��< ��<��<��<��<��<��<��<��<��<��<��<��< ��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<
��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��< ��<��<��<��<��<��<��<��<��<��<��<��<��<��< ��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   z�<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<
��<Z��<
��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��< ��<��<��<��<��<��< ��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<%��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<%��<��<`   `   ��<��<-��<��<��<2��<��<��<��<��<��<��<��<��<��<��<��<��<��<2��<��<��<-��<��<`   `   .��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<Y�<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   /��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<!��<��<��<��<��<��<��<��<��<��<��< ��<��<��<��<��<��<��<��<��<��<��<!��<`   `   ��<��<��<��<��<��< ��<��<��<��<��<��<��<��<��<��<��<��< ��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   
��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��< ��<��<��<��<��<��<��<��<��<��< ��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<z�<��<��<��<��<��<��<��<��<��<��<��<`   `   ǀ�<���<��<��<̀�<߀�<��<ـ�<��<ۀ�<Ӏ�<2��<��<2��<Ӏ�<ۀ�<��<ـ�<��<߀�<̀�<��<��<���<`   `   ���<ʀ�<���<؀�<���<ۀ�<	��<���<ހ�<Ā�<���<��<À�<��<���<Ā�<ހ�<���<	��<ۀ�<���<؀�<���<ʀ�<`   `   ���<��<���<���<܀�<���<��<���<ـ�<ڀ�<���<���<���<���<���<ڀ�<ـ�<���<��<���<܀�<���<���<��<`   `   ��<,��<��<���<��<̀�<���<Ѐ�<���<���<��<��<���<��<��<���<���<Ѐ�<���<̀�<��<���<��<,��<`   `   ��<���<���<���<���<���<Ѐ�<��<���<���<���<ۀ�<��<ۀ�<���<���<���<��<Ѐ�<���<���<���<���<���<`   `   ɀ�<؀�<܀�<���<��<΀�<���< ��<̀�<��< ��<���<��<���< ��<��<̀�< ��<���<΀�<��<���<܀�<؀�<`   `   Ҁ�<��<��<��<��<�<ڀ�<���<��<ހ�<���<܀�<���<܀�<���<ހ�<��<���<ڀ�<�<��<��<��<��<`   `   ܀�<ۀ�<��<Ҁ�<���<���<׀�<���<��<ۀ�<���<��<ǀ�<��<���<ۀ�<��<���<׀�<���<���<Ҁ�<��<ۀ�<`   `   ��<ۀ�<���<Հ�<���<��<؀�<Ā�<ۀ�<	��<Ӏ�<��< ��<��<Ӏ�<	��<ۀ�<Ā�<؀�<��<���<Հ�<���<ۀ�<`   `   ���<��<ƀ�<��<��<���<���<׀�<��<��<΀�<���<��<���<΀�<��<��<׀�<���<���<��<��<ƀ�<��<`   `   ��<���<��<π�<���<ڀ�<̀�<��<���<݀�<���<Ā�<���<Ā�<���<݀�<���<��<̀�<ڀ�<���<π�<��<���<`   `   ���< ��<���<À�<���<1��<��<؀�<���<π�<��<���<���<���<��<π�<���<؀�<��<1��<���<À�<���< ��<`   `   ǀ�<���<���<ۀ�<���<��<Հ�<؀�<��<��<��<��<��<��<��<��<��<؀�<Հ�<��<���<ۀ�<���<���<`   `   ��<��<��<��<��<���<��<��<Ā�<ـ�<���<Ѐ�<��<Ѐ�<���<ـ�<Ā�<��<��<���<��<��<��<��<`   `   ���<�<߀�<؀�<݀�<���<��<Ҁ�<���<ـ�<���<���<р�<���<���<ـ�<���<Ҁ�<��<���<݀�<؀�<߀�<�<`   `   ���<ˀ�<��<Ѐ�<��<ƀ�<���<ƀ�<��<���<р�<���<��<���<р�<���<��<ƀ�<���<ƀ�<��<Ѐ�<��<ˀ�<`   `   ���<р�<ڀ�<Հ�<��<ڀ�<�<"��<��<ˀ�<р�<��<Ҁ�<��<р�<ˀ�<��<"��<�<ڀ�<��<Հ�<ڀ�<р�<`   `   ـ�<Ҁ�<��<��<���<���<ƀ�<ހ�<ǀ�<���<���<ր�<���<ր�<���<���<ǀ�<ހ�<ƀ�<���<���<��<��<Ҁ�<`   `   ۀ�<�<���<��<Ѐ�<��<ǀ�<���<��<#��<��<���<
��<���<��<#��<��<���<ǀ�<��<Ѐ�<��<���<�<`   `   Ȁ�<���<��<Հ�<ـ�<���<��<��<��<��<���<���<��<���<���<��<��<��<��<���<ـ�<Հ�<��<���<`   `   π�<��<���<��<��<��<��<Ԁ�<Ѐ�<̀�<���<À�<���<À�<���<̀�<Ѐ�<Ԁ�<��<��<��<��<���<��<`   `   ڀ�<��<��<��<��<ـ�<��<ŀ�<Ӏ�<��<��<��<ʀ�<��<��<��<Ӏ�<ŀ�<��<ـ�<��<��<��<��<`   `   ��<��<���<���<Ā�<���<���<ր�<Ѐ�<���<���<��<���<��<���<���<Ѐ�<ր�<���<���<Ā�<���<���<��<`   `   ���<��<���<ۀ�<��<΀�<��<��<ˀ�<��<���<q��<���<q��<���<��<ˀ�<��<��<΀�<��<ۀ�<���<��<`   `   ��<2��<Ӏ�<ۀ�<��<ـ�<��<߀�<̀�<��<��<���<ǀ�<���<��<��<̀�<߀�<��<ـ�<��<ۀ�<Ӏ�<2��<`   `   À�<��<���<Ā�<ހ�<���<	��<ۀ�<���<؀�<���<ʀ�<���<ʀ�<���<؀�<���<ۀ�<	��<���<ހ�<Ā�<���<��<`   `   ���<���<���<ڀ�<ـ�<���<��<���<܀�<���<���<��<���<��<���<���<܀�<���<��<���<ـ�<ڀ�<���<���<`   `   ���<��<��<���<���<Ѐ�<���<̀�<��<���<��<,��<��<,��<��<���<��<̀�<���<Ѐ�<���<���<��<��<`   `   ��<ۀ�<���<���<���<��<Ѐ�<���<���<���<���<���<��<���<���<���<���<���<Ѐ�<��<���<���<���<ۀ�<`   `   ��<���< ��<��<̀�< ��<���<΀�<��<���<܀�<؀�<ɀ�<؀�<܀�<���<��<΀�<���< ��<̀�<��< ��<���<`   `   ���<܀�<���<ހ�<��<���<ڀ�<�<��<��<��<��<Ҁ�<��<��<��<��<�<ڀ�<���<��<ހ�<���<܀�<`   `   ǀ�<��<���<ۀ�<��<���<׀�<���<���<Ҁ�<��<ۀ�<܀�<ۀ�<��<Ҁ�<���<���<׀�<���<��<ۀ�<���<��<`   `    ��<��<Ӏ�<	��<ۀ�<Ā�<؀�<��<���<Հ�<���<ۀ�<��<ۀ�<���<Հ�<���<��<؀�<Ā�<ۀ�<	��<Ӏ�<��<`   `   ��<���<΀�<��<��<׀�<���<���<��<��<ƀ�<��<���<��<ƀ�<��<��<���<���<׀�<��<��<΀�<���<`   `   ���<Ā�<���<݀�<���<��<̀�<ڀ�<���<π�<��<���<��<���<��<π�<���<ڀ�<̀�<��<���<݀�<���<Ā�<`   `   ���<���<��<π�<���<؀�<��<1��<���<À�<���< ��<���< ��<���<À�<���<1��<��<؀�<���<π�<��<���<`   `   ��<��<��<��<��<؀�<Հ�<��<���<ۀ�<���<���<ǀ�<���<���<ۀ�<���<��<Հ�<؀�<��<��<��<��<`   `   ��<Ѐ�<���<ـ�<Ā�<��<��<���<��<��<��<��<��<��<��<��<��<���<��<��<Ā�<ـ�<���<Ѐ�<`   `   р�<���<���<ڀ�<���<Ҁ�<��<���<݀�<؀�<߀�<�<���<�<߀�<؀�<݀�<���<��<Ҁ�<���<ـ�<���<���<`   `   ��<���<р�<���<��<ƀ�<���<ƀ�<��<Ѐ�<��<ˀ�<���<ˀ�<��<Ѐ�<��<ƀ�<���<ƀ�<��<���<р�<���<`   `   Ҁ�<��<р�<ˀ�<��<"��<�<ڀ�<��<Հ�<ڀ�<р�<���<р�<ڀ�<Հ�<��<ڀ�<�<"��<��<ˀ�<р�<��<`   `   ���<ր�<���<���<ǀ�<ހ�<ƀ�<���<���<��<��<Ҁ�<ـ�<Ҁ�<��<��<���<���<ƀ�<ހ�<ǀ�<���<���<ր�<`   `   
��<���<��<#��<��<���<ǀ�<��<Ѐ�<��<���<�<ۀ�<�<���<��<Ѐ�<��<ǀ�<���<��<#��<��<���<`   `   ��<���<���<��<��<��<��<���<ـ�<Հ�<��<���<Ȁ�<���<��<Հ�<ـ�<���<��<��<��<��<���<���<`   `   ���<À�<���<̀�<Ѐ�<Ԁ�<��<��<��<��<���<��<π�<��<���<��<��<��<��<Ԁ�<Ѐ�<̀�<���<À�<`   `   ʀ�<��<��<��<Ӏ�<ŀ�<��<ـ�<��<��<��<��<ڀ�<��<��<��<��<ـ�<��<ŀ�<Ӏ�<��<��<��<`   `   ���<��<���<���<Ѐ�<ր�<���<���<Ā�<���<���<��<��<��<���<���<Ā�<���<���<ր�<Ѐ�<���<���<��<`   `   ���<q��<���<��<ˀ�<��<��<΀�<��<ۀ�<���<��<���<��<���<ۀ�<��<΀�<��<��<ˀ�<��<���<q��<`   `   ��<��<���<΁�<	��<ρ�<���<��<Ձ�<��<��<΁�<���<΁�<��<��<Ձ�<��<���<ρ�<	��<΁�<���<��<`   `   7��<0��<���<���<��<��<��<��<��<$��<���<Ё�<��<Ё�<���<$��<��<��<��<��<��<���<���<0��<`   `   ��<��<݁�<��<��<��<��<��<"��<��<��<���<5��<���<��<��<"��<��<��<��<��<��<݁�<��<`   `   ׁ�<���<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<���<`   `   ��<��<���<��<���<���<��<��<��<ˁ�<���<��<���<��<���<ˁ�<��<��<��<���<���<��<���<��<`   `   ��<��<ہ�<Ӂ�<��<؁�<��<݁�<	��<��<��<��<ځ�<��<��<��<	��<݁�<��<؁�<��<Ӂ�<ہ�<��<`   `   ��<���<݁�<ǁ�<���<��<��<�<?��<3��<���<6��<��<6��<���<3��<?��<�<��<��<���<ǁ�<݁�<���<`   `   Ɓ�<߁�<��<��<��<	��<%��<ف�<��<ށ�<Ɓ�<G��<���<G��<Ɓ�<ށ�<��<ف�<%��<	��<��<��<��<߁�<`   `   ��<���<$��<ρ�<��<��<��<%��<��<��<��<��<u��<��<��<��<��<%��<��<��<��<ρ�<$��<���<`   `   A��<��<��<ځ�<߁�<"��<��<$��<���<��<��<��<���<��<��<��<���<$��<��<"��<߁�<ځ�<��<��<`   `   ��<���<��<)��<ف�<��<Ё�<��<��<���<��< ��<7��< ��<��<���<��<��<Ё�<��<ف�<)��<��<���<`   `   ��<���<��<��<��<���<ځ�<��<��<��<��<Ӂ�<���<Ӂ�<��<��<��<��<ځ�<���<��<��<��<���<`   `   ��<��<Ӂ�<ԁ�<���<ځ�<���<���<��<���<��<��<'��<��<��<���<��<���<���<ځ�<���<ԁ�<Ӂ�<��<`   `   ��<��<��<��<��<���<Ձ�<��<܁�<��<���<���<D��<���<���<��<܁�<��<Ձ�<���<��<��<��<��<`   `   ��<ځ�<��<��<��<���<���<��<"��<1��<��<ԁ�<ہ�<ԁ�<��<1��<"��<��<���<���<��<��<��<ځ�<`   `   +��<��< ��<��<��<���<��<���<��<��<��<��<��<��<��<��<��<���<��<���<��<��< ��<��<`   `   "��<	��<��<���<��<��<2��<с�<́�<���<؁�<��<��<��<؁�<���<́�<с�<2��<��<��<���<��<	��<`   `   ��<��<���<��<���<߁�<+��<���<��<��<��<��<܁�<��<��<��<��<���<+��<߁�<���<��<���<��<`   `   ��<��<���<)��<���<���<܁�<���<��<́�<ف�<��<��<��<ف�<́�<��<���<܁�<���<���<)��<���<��<`   `   ��<��<��<��<��<��<��<���<��<���<��<��<��<��<��<���<��<���<��<��<��<��<��<��<`   `   ���<��<���<���<́�<��<!��<܁�<���<���<��<%��<��<%��<��<���<���<܁�<!��<��<́�<���<���<��<`   `   Ɂ�<���<��<��<���<ځ�<��<΁�<%��<��<Ɂ�<���<߁�<���<Ɂ�<��<%��<΁�<��<ځ�<���<��<��<���<`   `   ʁ�<��<��<%��<��<��<���<���<��<ށ�<ȁ�<���<0��<���<ȁ�<ށ�<��<���<���<��<��<%��<��<��<`   `   Ё�<��<��<��<ʁ�< ��<��<��<���<ȁ�<���<(��<E��<(��<���<ȁ�<���<��<��< ��<ʁ�<��<��<��<`   `   ���<΁�<��<��<Ձ�<��<���<ρ�<	��<΁�<���<��<��<��<���<΁�<	��<ρ�<���<��<Ձ�<��<��<΁�<`   `   ��<Ё�<���<$��<��<��<��<��<��<���<���<0��<7��<0��<���<���<��<��<��<��<��<$��<���<Ё�<`   `   5��<���<��<��<"��<��<��<��<��<��<݁�<��<��<��<݁�<��<��<��<��<��<"��<��<��<���<`   `   ��<��<��<��<��<��<��<��<��<��<��<���<ׁ�<���<��<��<��<��<��<��<��<��<��<��<`   `   ���<��<���<ˁ�<��<��<��<���<���<��<���<��<��<��<���<��<���<���<��<��<��<ˁ�<���<��<`   `   ځ�<��<��<��<	��<݁�<��<؁�<��<Ӂ�<ہ�<��<��<��<ہ�<Ӂ�<��<؁�<��<݁�<	��<��<��<��<`   `   ��<6��<���<3��<?��<�<��<��<���<ǁ�<݁�<���<��<���<݁�<ǁ�<���<��<��<�<?��<3��<���<6��<`   `   ���<G��<Ɓ�<ށ�<��<ف�<%��<	��<��<��<��<߁�<Ɓ�<߁�<��<��<��<	��<%��<ف�<��<ށ�<Ɓ�<G��<`   `   u��<��<��<��<��<%��<��<��<��<ρ�<$��<���<��<���<$��<ρ�<��<��<��<%��<��<��<��<��<`   `   ���<��<��<��<���<$��<��<"��<߁�<ځ�<��<��<A��<��<��<ځ�<߁�<"��<��<$��<���<��<��<��<`   `   7��< ��<��<���<��<��<Ё�<��<ف�<)��<��<���<��<���<��<)��<ف�<��<Ё�<��<��<���<��< ��<`   `   ���<Ӂ�<��<��<��<��<ځ�<���<��<��<��<���<��<���<��<��<��<���<ځ�<��<��<��<��<Ӂ�<`   `   '��<��<��<���<��<���<���<ځ�<���<ԁ�<Ӂ�<��<��<��<Ӂ�<ԁ�<���<ځ�<���<���<��<���<��<��<`   `   D��<���<���<��<܁�<��<Ձ�<���<��<��<��<��<��<��<��<��<��<���<Ձ�<��<܁�<��<���<���<`   `   ہ�<ԁ�<��<1��<"��<��<���<���<��<��<��<ځ�<��<ځ�<��<��<��<���<���<��<"��<1��<��<ԁ�<`   `   ��<��<��<��<��<���<��<���<��<��< ��<��<+��<��< ��<��<��<���<��<���<��<��<��<��<`   `   ��<��<؁�<���<́�<с�<2��<��<��<���<��<	��<"��<	��<��<���<��<��<2��<с�<́�<���<؁�<��<`   `   ܁�<��<��<��<��<���<+��<߁�<���<��<���<��<��<��<���<��<���<߁�<+��<���<��<��<��<��<`   `   ��<��<ف�<́�<��<���<܁�<���<���<)��<���<��<��<��<���<)��<���<���<܁�<���<��<́�<ف�<��<`   `   ��<��<��<���<��<���<��<��<��<��<��<��<��<��<��<��<��<��<��<���<��<���<��<��<`   `   ��<%��<��<���<���<܁�<!��<��<́�<���<���<��<���<��<���<���<́�<��<!��<܁�<���<���<��<%��<`   `   ߁�<���<Ɂ�<��<%��<΁�<��<ځ�<���<��<��<���<Ɂ�<���<��<��<���<ځ�<��<΁�<%��<��<Ɂ�<���<`   `   0��<���<ȁ�<ށ�<��<���<���<��<��<%��<��<��<ʁ�<��<��<%��<��<��<���<���<��<ށ�<ȁ�<���<`   `   E��<(��<���<ȁ�<���<��<��< ��<ʁ�<��<��<��<Ё�<��<��<��<ʁ�< ��<��<��<���<ȁ�<���<(��<`   `   ���<���<��<��<:��<A��<��<B��<��<#��<��<��<{��<��<��<#��<��<B��<��<A��<:��<��<��<���<`   `   ���<��<���<$��<(��<��<-��<B��<��<��<-��<&��<m��<&��<-��<��<��<B��<-��<��<(��<$��<���<��<`   `   Q��<��<��<T��<��<���<��<��<҂�<ǂ�<#��<��<��<��<#��<ǂ�<҂�<��<��<���<��<T��<��<��<`   `   \��<��<��<-��<߂�<;��<��<��<@��<-��<��<��<��<��<��<-��<@��<��<��<;��<߂�<-��<��<��<`   `   ��< ��<Q��< ��<��<T��<��<��<D��<?��<��<3��<o��<3��<��<?��<D��<��<��<T��<��< ��<Q��< ��<`   `   ��<��<C��<��<��<��<���<��<��<���<��<��<��<��<��<���<��<��<���<��<��<��<C��<��<`   `   D��<��<��<��<<��<��<<��<M��<���<��<+��<��<܂�<��<+��<��<���<M��<<��<��<<��<��<��<��<`   `   X��<��<$��<&��<<��<߂�<��<K��<��<2��<3��<>��<��<>��<3��<2��<��<K��<��<߂�<<��<&��<$��<��<`   `   ��<��<6��<��<��<���<ł�<��<���<%��<��<��<��<��<��<%��<���<��<ł�<���<��<��<6��<��<`   `   ��<��<%��<��<(��<&��< ��<��<��<6��<��<��<��<��<��<6��<��<��< ��<&��<(��<��<%��<��<`   `   7��<��<��<��<%��<$��<3��<���<��<U��<��<��<1��<��<��<U��<��<���<3��<$��<%��<��<��<��<`   `   W��<H��<��</��<��<��<9��<(��<��<>��<��<��<3��<��<��<>��<��<(��<9��<��<��</��<��<H��<`   `   ��<-��<��<4��<<��<2��<a��<@��<��<	��<��<��<%��<��<��<	��<��<@��<a��<2��<<��<4��<��<-��<`   `   ���<&��<#��<��<)��<A��<��<
��<!��<��<.��<��<��<��<.��<��<!��<
��<��<A��<)��<��<#��<&��<`   `   2��<,��<���<���<��<*��<��<*��<'��<˂�<A��<F��<���<F��<A��<˂�<'��<*��<��<*��<��<���<���<,��<`   `   ��<��<��<��<$��<)��<8��<D��<��<���<��<!��<Ղ�<!��<��<���<��<D��<8��<)��<$��<��<��<��<`   `   ۂ�<��<3��<&��<#��<��<��<���<��<3��< ��<��<��<��< ��<3��<��<���<��<��<#��<&��<3��<��<`   `   ��<5��<)��<��<7��<*��<��<��<;��<X��<-��<I��<k��<I��<-��<X��<;��<��<��<*��<7��<��<)��<5��<`   `   ��<(��< ��<���<U��<;��<��<;��<'��<��<��<��<��<��<��<��<'��<;��<��<;��<U��<���< ��<(��<`   `   ��<��<��<:��<L��<��<��<��<��<+��<;��<���<��<���<;��<+��<��<��<��<��<L��<:��<��<��<`   `   ���<��<��<D��<'��<���<��<&��<��<7��<>��</��<Z��</��<>��<7��<��<&��<��<���<'��<D��<��<��<`   `   ?��<(��<��< ��<��<��<$��<A��<��<���< ��<��<$��<��< ��<���<��<A��<$��<��<��< ��<��<(��<`   `   L��<1��<&��<��<��<=��<��<��<���<��<V��<���<��<���<V��<��<���<��<��<=��<��<��<&��<1��<`   `   S��<��<��<��<��<E��<
��<)��< ��<)��<v��<"��<ӂ�<"��<v��<)��< ��<)��<
��<E��<��<��<��<��<`   `   {��<��<��<#��<��<B��<��<A��<:��<��<��<���<���<���<��<��<:��<A��<��<B��<��<#��<��<��<`   `   m��<&��<-��<��<��<B��<-��<��<(��<$��<���<��<���<��<���<$��<(��<��<-��<B��<��<��<-��<&��<`   `   ��<��<#��<ǂ�<҂�<��<��<���<��<T��<��<��<Q��<��<��<T��<��<���<��<��<҂�<ǂ�<#��<��<`   `   ��<��<��<-��<@��<��<��<;��<߂�<-��<��<��<\��<��<��<-��<߂�<;��<��<��<@��<-��<��<��<`   `   o��<3��<��<?��<D��<��<��<T��<��< ��<Q��< ��<��< ��<Q��< ��<��<T��<��<��<D��<?��<��<3��<`   `   ��<��<��<���<��<��<���<��<��<��<C��<��<��<��<C��<��<��<��<���<��<��<���<��<��<`   `   ܂�<��<+��<��<���<M��<<��<��<<��<��<��<��<D��<��<��<��<<��<��<<��<M��<���<��<+��<��<`   `   ��<>��<3��<2��<��<K��<��<߂�<<��<&��<$��<��<X��<��<$��<&��<<��<߂�<��<K��<��<2��<3��<>��<`   `   ��<��<��<%��<���<��<ł�<���<��<��<6��<��<��<��<6��<��<��<���<ł�<��<���<%��<��<��<`   `   ��<��<��<6��<��<��< ��<&��<(��<��<%��<��<��<��<%��<��<(��<&��< ��<��<��<6��<��<��<`   `   1��<��<��<U��<��<���<3��<$��<%��<��<��<��<7��<��<��<��<%��<$��<3��<���<��<U��<��<��<`   `   3��<��<��<>��<��<(��<9��<��<��</��<��<H��<W��<H��<��</��<��<��<9��<(��<��<>��<��<��<`   `   %��<��<��<	��<��<@��<a��<2��<<��<4��<��<-��<��<-��<��<4��<<��<2��<a��<@��<��<	��<��<��<`   `   ��<��<.��<��<!��<
��<��<A��<)��<��<#��<&��<���<&��<#��<��<)��<A��<��<
��<!��<��<.��<��<`   `   ���<F��<A��<˂�<'��<*��<��<*��<��<���<���<,��<2��<,��<���<���<��<*��<��<*��<'��<˂�<A��<F��<`   `   Ղ�<!��<��<���<��<D��<8��<)��<$��<��<��<��<��<��<��<��<$��<)��<8��<D��<��<���<��<!��<`   `   ��<��< ��<3��<��<���<��<��<#��<&��<3��<��<ۂ�<��<3��<&��<#��<��<��<���<��<3��< ��<��<`   `   k��<I��<-��<X��<;��<��<��<*��<7��<��<)��<5��<��<5��<)��<��<7��<*��<��<��<;��<X��<-��<I��<`   `   ��<��<��<��<'��<;��<��<;��<U��<���< ��<(��<��<(��< ��<���<U��<;��<��<;��<'��<��<��<��<`   `   ��<���<;��<+��<��<��<��<��<L��<:��<��<��<��<��<��<:��<L��<��<��<��<��<+��<;��<���<`   `   Z��</��<>��<7��<��<&��<��<���<'��<D��<��<��<���<��<��<D��<'��<���<��<&��<��<7��<>��</��<`   `   $��<��< ��<���<��<A��<$��<��<��< ��<��<(��<?��<(��<��< ��<��<��<$��<A��<��<���< ��<��<`   `   ��<���<V��<��<���<��<��<=��<��<��<&��<1��<L��<1��<&��<��<��<=��<��<��<���<��<V��<���<`   `   ӂ�<"��<v��<)��< ��<)��<
��<E��<��<��<��<��<S��<��<��<��<��<E��<
��<)��< ��<)��<v��<"��<`   `   ���<w��<K��<u��<��<N��<\��<��<s��<_��<4��<<��<G��<<��<4��<_��<s��<��<\��<N��<��<u��<K��<w��<`   `   @��<���<���<O��<#��<P��<=��<-��<���<v��<\��<C��<��<C��<\��<v��<���<-��<=��<P��<#��<O��<���<���<`   `   ��<]��<`��<;��<l��<Z��<G��<^��<|��<c��<q��<U��<��<U��<q��<c��<|��<^��<G��<Z��<l��<;��<`��<]��<`   `   .��<g��<4��<-��<y��<G��<Q��<O��<0��<>��<G��<Q��<Z��<Q��<G��<>��<0��<O��<Q��<G��<y��<-��<4��<g��<`   `   c��<Y��<��<&��<^��<9��<O��<r��<L��<L��<G��<@��<`��<@��<G��<L��<L��<r��<O��<9��<^��<&��<��<Y��<`   `   J��<<��<C��<]��<W��<D��<C��<���<f��<D��<w��<@��<V��<@��<w��<D��<f��<���<C��<D��<W��<]��<C��<<��<`   `   I��<E��<n��<Z��<2��<\��<!��<c��<5��<D��<x��<+��<s��<+��<x��<D��<5��<c��<!��<\��<2��<Z��<n��<E��<`   `   ]��<@��<<��<'��<0��<���<M��<7��<K��<j��<,��<���<���<���<,��<j��<K��<7��<M��<���<0��<'��<<��<@��<`   `   h��<R��<9��<K��<Z��<���<{��<D��<a��<d��<-��<L��<���<L��<-��<d��<a��<D��<{��<���<Z��<K��<9��<R��<`   `   W��<��<W��<X��<g��<E��<r��<R��<S��<O��<\��<q��<F��<q��<\��<O��<S��<R��<r��<E��<g��<X��<W��<��<`   `   ��<u��<A��<��<f��<)��<Z��<V��<c��<V��<L��<C��<��<C��<L��<V��<c��<V��<Z��<)��<f��<��<A��<u��<`   `   ��<[��<J��<#��<c��</��<2��<��<?��<?��<P��<���<S��<���<P��<?��<?��<��<2��</��<c��<#��<J��<[��<`   `   ��<J��<I��<I��<C��<C��<U��<+��<P��<H��<X��<k��<G��<k��<X��<H��<P��<+��<U��<C��<C��<I��<I��<J��<`   `   N��<Y��<@��<W��<#��</��<T��<;��<���<t��<F��<.��<0��<.��<F��<t��<���<;��<T��</��<#��<W��<@��<Y��<`   `   H��<j��<`��<y��<M��<>��<?��<��<S��<k��<<��<I��<���<I��<<��<k��<S��<��<?��<>��<M��<y��<`��<j��<`   `   3��<X��<Z��<c��<Z��<Y��<\��<R��<m��<���<\��<H��<���<H��<\��<���<m��<R��<\��<Y��<Z��<c��<Z��<X��<`   `   S��<O��<M��<P��<F��<'��<"��<g��<w��<d��<S��<8��<B��<8��<S��<d��<w��<g��<"��<'��<F��<P��<M��<O��<`   `   M��<I��<Z��<[��<b��<G��<*��<L��<��<��<+��<3��<0��<3��<+��<��<��<L��<*��<G��<b��<[��<Z��<I��<`   `   J��<W��<[��<��< ��<]��<j��<S��<(��<N��<i��<X��<d��<X��<i��<N��<(��<S��<j��<]��< ��<��<[��<W��<`   `   h��<c��<d��<.��<��<G��<W��<H��<X��<|��<H��<4��<|��<4��<H��<|��<X��<H��<W��<G��<��<.��<d��<c��<`   `   }��<T��<Y��<j��<V��<}��<Z��<Q��<G��<6��<��<��<\��<��<��<6��<G��<Q��<Z��<}��<V��<j��<Y��<T��<`   `   T��<B��<=��<3��<H��<n��<L��<^��<>��<L��<���<j��<|��<j��<���<L��<>��<^��<L��<n��<H��<3��<=��<B��<`   `   ��<9��<X��<,��<8��<7��<1��<M��<F��<e��<N��<Q��<���<Q��<N��<e��<F��<M��<1��<7��<8��<,��<X��<9��<`   `   *��<@��<X��<Z��<_��<'��<U��<L��<=��<h��<��<'��<���<'��<��<h��<=��<L��<U��<'��<_��<Z��<X��<@��<`   `   G��<<��<4��<_��<s��<��<\��<N��<��<u��<K��<w��<���<w��<K��<u��<��<N��<\��<��<s��<_��<4��<<��<`   `   ��<C��<\��<v��<���<-��<=��<P��<#��<O��<���<���<@��<���<���<O��<#��<P��<=��<-��<���<v��<\��<C��<`   `   ��<U��<q��<c��<|��<^��<G��<Z��<l��<;��<`��<]��<��<]��<`��<;��<l��<Z��<G��<^��<|��<c��<q��<U��<`   `   Z��<Q��<G��<>��<0��<O��<Q��<G��<y��<-��<4��<g��<.��<g��<4��<-��<y��<G��<Q��<O��<0��<>��<G��<Q��<`   `   `��<@��<G��<L��<L��<r��<O��<9��<^��<&��<��<Y��<c��<Y��<��<&��<^��<9��<O��<r��<L��<L��<G��<@��<`   `   V��<@��<w��<D��<f��<���<C��<D��<W��<]��<C��<<��<J��<<��<C��<]��<W��<D��<C��<���<f��<D��<w��<@��<`   `   s��<+��<x��<D��<5��<c��<!��<\��<2��<Z��<n��<E��<I��<E��<n��<Z��<2��<\��<!��<c��<5��<D��<x��<+��<`   `   ���<���<,��<j��<K��<7��<M��<���<0��<'��<<��<@��<]��<@��<<��<'��<0��<���<M��<7��<K��<j��<,��<���<`   `   ���<L��<-��<d��<a��<D��<{��<���<Z��<K��<9��<R��<h��<R��<9��<K��<Z��<���<{��<D��<a��<d��<-��<L��<`   `   F��<q��<\��<O��<S��<R��<r��<E��<g��<X��<W��<��<W��<��<W��<X��<g��<E��<r��<R��<S��<O��<\��<q��<`   `   ��<C��<L��<V��<c��<V��<Z��<)��<f��<��<A��<u��<��<u��<A��<��<f��<)��<Z��<V��<c��<V��<L��<C��<`   `   S��<���<P��<?��<?��<��<2��</��<c��<#��<J��<[��<��<[��<J��<#��<c��</��<2��<��<?��<?��<P��<���<`   `   G��<k��<X��<H��<P��<+��<U��<C��<C��<I��<I��<J��<��<J��<I��<I��<C��<C��<U��<+��<P��<H��<X��<k��<`   `   0��<.��<F��<t��<���<;��<T��</��<#��<W��<@��<Y��<N��<Y��<@��<W��<#��</��<T��<;��<���<t��<F��<.��<`   `   ���<I��<<��<k��<S��<��<?��<>��<M��<y��<`��<j��<H��<j��<`��<y��<M��<>��<?��<��<S��<k��<<��<I��<`   `   ���<H��<\��<���<m��<R��<\��<Y��<Z��<c��<Z��<X��<3��<X��<Z��<c��<Z��<Y��<\��<R��<m��<���<\��<H��<`   `   B��<8��<S��<d��<w��<g��<"��<'��<F��<P��<M��<O��<S��<O��<M��<P��<F��<'��<"��<g��<w��<d��<S��<8��<`   `   0��<3��<+��<��<��<L��<*��<G��<b��<[��<Z��<I��<M��<I��<Z��<[��<b��<G��<*��<L��<��<��<+��<3��<`   `   d��<X��<i��<N��<(��<S��<j��<]��< ��<��<[��<W��<J��<W��<[��<��< ��<]��<j��<S��<(��<N��<i��<X��<`   `   |��<4��<H��<|��<X��<H��<W��<G��<��<.��<d��<c��<h��<c��<d��<.��<��<G��<W��<H��<X��<|��<H��<4��<`   `   \��<��<��<6��<G��<Q��<Z��<}��<V��<j��<Y��<T��<}��<T��<Y��<j��<V��<}��<Z��<Q��<G��<6��<��<��<`   `   |��<j��<���<L��<>��<^��<L��<n��<H��<3��<=��<B��<T��<B��<=��<3��<H��<n��<L��<^��<>��<L��<���<j��<`   `   ���<Q��<N��<e��<F��<M��<1��<7��<8��<,��<X��<9��<��<9��<X��<,��<8��<7��<1��<M��<F��<e��<N��<Q��<`   `   ���<'��<��<h��<=��<L��<U��<'��<_��<Z��<X��<@��<*��<@��<X��<Z��<_��<'��<U��<L��<=��<h��<��<'��<`   `   k��<���<���<ʅ�<���<u��<���<���<g��<C��<���<���<u��<���<���<C��<g��<���<���<u��<���<ʅ�<���<���<`   `   ���<b��<S��<s��<���<���<���<l��<p��<Z��<t��<���<|��<���<t��<Z��<p��<l��<���<���<���<s��<S��<b��<`   `   ���<���<p��<Z��<���<���<���<���<���<���<d��<���<ƅ�<���<d��<���<���<���<���<���<���<Z��<p��<���<`   `   W��<���<���<���<���<I��<���<���<h��<���<��<���<���<���<��<���<h��<���<���<I��<���<���<���<���<`   `   u��<���<���<���<���<_��<���<[��<`��<���<���<|��<9��<|��<���<���<`��<[��<���<_��<���<���<���<���<`   `   ���<���<m��<���<���<���<���<i��<���<���<���<���<���<���<���<���<���<i��<���<���<���<���<m��<���<`   `   t��<���<���<���<e��<���<`��<^��<���<k��<���<���<��<���<���<k��<���<^��<`��<���<e��<���<���<���<`   `   O��<���<���<���<d��<���<���<���<���<k��<���<l��<���<l��<���<k��<���<���<���<���<d��<���<���<���<`   `   d��<���<{��<���<e��<���<���<���<���<b��<Ņ�<~��<?��<~��<Ņ�<b��<���<���<���<���<e��<���<{��<���<`   `   v��<���<v��<���<b��<B��<`��<]��<��<K��<���<���<m��<���<���<K��<��<]��<`��<B��<b��<���<v��<���<`   `   ���<|��<���<���<���<���<���<���<���<a��<v��<���<���<���<v��<a��<���<���<���<���<���<���<���<|��<`   `   ą�<���<���<���<���<ȅ�<���<���<���<���<r��<���<���<���<r��<���<���<���<���<ȅ�<���<���<���<���<`   `   ��<���<���<���<���<���<k��<���<���<���<���<���<f��<���<���<���<���<���<k��<���<���<���<���<���<`   `   ���<���<a��<���<���<���<���<���<}��<i��<���<���<���<���<���<i��<}��<���<���<���<���<���<a��<���<`   `   X��<{��<y��<���<���<���<���<���<_��<���<y��<e��<���<e��<y��<���<_��<���<���<���<���<���<y��<{��<`   `   ���<���<���<w��<x��<���<���<m��<U��<���<���<Z��<���<Z��<���<���<U��<m��<���<���<x��<w��<���<���<`   `   ���<���<l��<l��<n��<Å�<���<���<p��<k��<���<�<ȅ�<�<���<k��<p��<���<���<Å�<n��<l��<l��<���<`   `   ���<a��<y��<���<���<���<���<���<���<���<���<���<b��<���<���<���<���<���<���<���<���<���<y��<a��<`   `   ���<s��<���<؅�<���<x��<���<���<���<���<���<���<p��<���<���<���<���<���<���<x��<���<؅�<���<s��<`   `   ���<{��<q��<���<���<���<���<���<���<j��<���<ą�<Ņ�<ą�<���<j��<���<���<���<���<���<���<q��<{��<`   `   ���<v��<p��<���<���<���<u��<���<���<l��<���<���<Z��<���<���<l��<���<���<u��<���<���<���<p��<v��<`   `   ���<���<���<���<���<~��<m��<u��<���<���<���<���<<��<���<���<���<���<u��<m��<~��<���<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<l��<c��<���<S��<���<c��<l��<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<���<���<���<~��<���<���<g��<���<h��<���<g��<���<���<~��<���<���<���<���<���<���<`   `   u��<���<���<C��<g��<���<���<u��<���<ʅ�<���<���<k��<���<���<ʅ�<���<u��<���<���<g��<C��<���<���<`   `   |��<���<t��<Z��<p��<l��<���<���<���<s��<S��<b��<���<b��<S��<s��<���<���<���<l��<p��<Z��<t��<���<`   `   ƅ�<���<d��<���<���<���<���<���<���<Z��<p��<���<���<���<p��<Z��<���<���<���<���<���<���<d��<���<`   `   ���<���<��<���<h��<���<���<I��<���<���<���<���<W��<���<���<���<���<I��<���<���<h��<���<��<���<`   `   9��<|��<���<���<`��<[��<���<_��<���<���<���<���<u��<���<���<���<���<_��<���<[��<`��<���<���<|��<`   `   ���<���<���<���<���<i��<���<���<���<���<m��<���<���<���<m��<���<���<���<���<i��<���<���<���<���<`   `   ��<���<���<k��<���<^��<`��<���<e��<���<���<���<t��<���<���<���<e��<���<`��<^��<���<k��<���<���<`   `   ���<l��<���<k��<���<���<���<���<d��<���<���<���<O��<���<���<���<d��<���<���<���<���<k��<���<l��<`   `   ?��<~��<Ņ�<b��<���<���<���<���<e��<���<{��<���<d��<���<{��<���<e��<���<���<���<���<b��<Ņ�<~��<`   `   m��<���<���<K��<��<]��<`��<B��<b��<���<v��<���<v��<���<v��<���<b��<B��<`��<]��<��<K��<���<���<`   `   ���<���<v��<a��<���<���<���<���<���<���<���<|��<���<|��<���<���<���<���<���<���<���<a��<v��<���<`   `   ���<���<r��<���<���<���<���<ȅ�<���<���<���<���<ą�<���<���<���<���<ȅ�<���<���<���<���<r��<���<`   `   f��<���<���<���<���<���<k��<���<���<���<���<���<��<���<���<���<���<���<k��<���<���<���<���<���<`   `   ���<���<���<i��<}��<���<���<���<���<���<a��<���<���<���<a��<���<���<���<���<���<}��<i��<���<���<`   `   ���<e��<y��<���<_��<���<���<���<���<���<y��<{��<X��<{��<y��<���<���<���<���<���<_��<���<y��<e��<`   `   ���<Z��<���<���<U��<m��<���<���<x��<w��<���<���<���<���<���<w��<x��<���<���<m��<U��<���<���<Z��<`   `   ȅ�<�<���<k��<p��<���<���<Å�<n��<l��<l��<���<���<���<l��<l��<n��<Å�<���<���<p��<k��<���<�<`   `   b��<���<���<���<���<���<���<���<���<���<y��<a��<���<a��<y��<���<���<���<���<���<���<���<���<���<`   `   p��<���<���<���<���<���<���<x��<���<؅�<���<s��<���<s��<���<؅�<���<x��<���<���<���<���<���<���<`   `   Ņ�<ą�<���<j��<���<���<���<���<���<���<q��<{��<���<{��<q��<���<���<���<���<���<���<j��<���<ą�<`   `   Z��<���<���<l��<���<���<u��<���<���<���<p��<v��<���<v��<p��<���<���<���<u��<���<���<l��<���<���<`   `   <��<���<���<���<���<u��<m��<~��<���<���<���<���<���<���<���<���<���<~��<m��<u��<���<���<���<���<`   `   S��<���<c��<l��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<l��<c��<���<`   `   h��<���<g��<���<���<~��<���<���<���<���<���<���<���<���<���<���<���<���<���<~��<���<���<g��<���<`   `   ���<߆�<��<���<��<Ն�<Ɇ�<$��<��<��<��<�<ц�<�<��<��<��<$��<Ɇ�<Ն�<��<���<��<߆�<`   `   ��<���<��<���<݆�<׆�<ֆ�<	��<͆�<��<���<Ά�<��<Ά�<���<��<͆�<	��<ֆ�<׆�<݆�<���<��<���<`   `   `��<Ն�<��<��<���<Ɇ�<�<ņ�<���<��<���<���<Ɔ�<���<���<��<���<ņ�<�<Ɇ�<���<��<��<Ն�<`   `   ���<���<Ԇ�<���<���<���<���<���<���<���<ˆ�<߆�<���<߆�<ˆ�<���<���<���<���<���<���<���<Ԇ�<���<`   `   ֆ�<ņ�<��<�<ǆ�<��<ֆ�<Ć�<��<��<���<8��<���<8��<���<��<��<Ć�<ֆ�<��<Ȇ�<�<��<ņ�<`   `   ���<��<݆�<ֆ�<Ɔ�<��<���<���<���<φ�<���<��<Ն�<��<���<φ�<���<���<���<��<Ɔ�<ֆ�<݆�<��<`   `   ���<��<���<��<��<͆�<��<���<��<ц�<׆�<���<���<���<׆�<ц�<��<���<��<͆�<��<��<���<��<`   `   ݆�<��<���<���<��<���<��<���<̆�<���<��<��<��<��<��<���<̆�<���<��<���<��<���<���<��<`   `   Ɇ�<	��<���<ц�<���<��<��<Ն�<��<Ć�<͆�<І�< ��<І�<͆�<Ć�<��<Ն�<��<��<���<ц�<���<	��<`   `   ׆�<��<ц�<ǆ�<��<#��<��<ņ�<	��<��<���<���<���<���<���<��<	��<ņ�<��<#��<��<ǆ�<ц�<��<`   `   !��<φ�<��<Ԇ�<�<���<چ�<φ�<���<&��<��<���<��<���<��<&��<���<φ�<چ�<���<�<Ԇ�<��<φ�<`   `   ��<���<߆�<���<���<Ɇ�<Ɔ�<��<���<��<���<���<��<���<���<��<���<��<Ɔ�<Ɇ�<���<���<߆�<���<`   `   ���<���<���<׆�<���<��<���<܆�<ц�<��<؆�<���<Ɇ�<���<؆�<��<ц�<܆�<���<��<���<׆�<���<���<`   `   ���<��<��<ֆ�<���<��<���<Ɇ�<ʆ�<Ć�<��<���<ن�<���<��<Ć�<ʆ�<Ɇ�<���<��<���<ֆ�<��<��<`   `   ��<��<��<���<��<���<���<���<��<��<��<��<Ȇ�<��<��<��<��<���<���<���<��<���<��<��<`   `   �<І�<��<��<���<���<���< ��<��<φ�<܆�<ӆ�<���<ӆ�<܆�<φ�<��< ��<���<���<���<��<��<І�<`   `   ���<���<��<��<���<��<���<ǆ�<��<���<ˆ�<��<ц�<��<ˆ�<���<��<ǆ�<���<��<���<��<��<���<`   `   ���<��<���<���<���<φ�<͆�<���<���<��<ц�<��<��<��<ц�<��<���<���<͆�<φ�<���<���<���<��<`   `   ؆�<��<ӆ�<���<܆�<Ɇ�<Ն�<���<Ć�<چ�<���<���<ǆ�<���<���<چ�<Ć�<���<Ն�<Ɇ�<܆�<���<ӆ�<��<`   `   Ԇ�<��<ц�<ʆ�<
��<���<��<��<ˆ�<���<ۆ�<ӆ�<���<ӆ�<ۆ�<���<ˆ�<��<��<���<
��<ʆ�<ц�<��<`   `   ���<���<���<Ԇ�<ӆ�<Ȇ�<��<��<��<���<���<��<؆�<��<���<���<��<��<��<Ȇ�<ӆ�<Ԇ�<���<���<`   `   ؆�<��<��<܆�<͆�<ކ�<��<ǆ�<���<ކ�<���<҆�<+��<҆�<���<ކ�<���<ǆ�<��<ކ�<͆�<܆�<��<��<`   `   ���<���<���<Ć�<ǆ�<ʆ�<���<؆�<ˆ�<ӆ�<ن�<��<ن�<��<ن�<ӆ�<ˆ�<؆�<���<ʆ�<ǆ�<Ć�<���<���<`   `   ��<���<���<܆�<Ć�<���<���<Æ�<��<���<8��<3��<���<3��<8��<���<��<Æ�<���<���<Ć�<܆�<���<���<`   `   ц�<�<��<��<��<$��<Ɇ�<Ն�<��<���<��<߆�<���<߆�<��<���<��<Ն�<Ɇ�<$��<��<��<��<�<`   `   ��<Ά�<���<��<͆�<	��<ֆ�<׆�<݆�<���<��<���<��<���<��<���<݆�<׆�<ֆ�<	��<͆�<��<���<Ά�<`   `   Ɔ�<���<���<��<���<ņ�<�<Ɇ�<���<��<��<Ն�<`��<Ն�<��<��<���<Ɇ�<�<ņ�<���<��<���<���<`   `   ���<߆�<ˆ�<���<���<���<���<���<���<���<Ԇ�<���<���<���<Ԇ�<���<���<���<���<���<���<���<ˆ�<߆�<`   `   ���<8��<���<��<��<Ć�<ֆ�<��<ǆ�<�<��<ņ�<ֆ�<ņ�<��<�<ǆ�<��<ֆ�<Ć�<��<��<���<8��<`   `   Ն�<��<���<φ�<���<���<���<��<Ɔ�<ֆ�<݆�<��<���<��<݆�<ֆ�<Ɔ�<��<���<���<���<φ�<���<��<`   `   ���<���<׆�<ц�<��<���<��<͆�<��<��<���<��<���<��<���<��<��<͆�<��<���<��<ц�<׆�<���<`   `   ��<��<��<���<̆�<���<��<���<��<���<���<��<݆�<��<���<���<��<���<��<���<̆�<���<��<��<`   `    ��<І�<͆�<Ć�<��<Ն�<��<��<���<ц�<���<	��<Ɇ�<	��<���<ц�<���<��<��<Ն�<��<Ć�<͆�<І�<`   `   ���<���<���<��<	��<ņ�<��<#��<��<ǆ�<ц�<��<׆�<��<ц�<ǆ�<��<#��<��<ņ�<	��<��<���<���<`   `   ��<���<��<&��<���<φ�<چ�<���<�<Ԇ�<��<φ�<!��<φ�<��<Ԇ�<�<���<چ�<φ�<���<&��<��<���<`   `   ��<���<���<��<���<��<Ɔ�<Ɇ�<���<���<߆�<���<��<���<߆�<���<���<Ɇ�<Ɔ�<��<���<��<���<���<`   `   Ɇ�<���<؆�<��<ц�<܆�<���<��<���<׆�<���<���<���<���<���<׆�<���<��<���<܆�<ц�<��<؆�<���<`   `   ن�<���<��<Ć�<ʆ�<Ɇ�<���<��<���<ֆ�<��<��<���<��<��<ֆ�<���<��<���<Ɇ�<ʆ�<Ć�<��<���<`   `   Ȇ�<��<��<��<��<���<���<���<��<���<��<��<��<��<��<���<��<���<���<���<��<��<��<��<`   `   ���<ӆ�<܆�<φ�<��< ��<���<���<���<��<��<І�<�<І�<��<��<���<���<���< ��<��<φ�<܆�<ӆ�<`   `   ц�<��<ˆ�<���<��<ǆ�<���<��<���<��<��<���<���<���<��<��<���<��<���<ǆ�<��<���<ˆ�<��<`   `   ��<��<ц�<��<���<���<͆�<φ�<���<���<���<��<���<��<���<���<���<φ�<͆�<���<���<��<ц�<��<`   `   ǆ�<���<���<چ�<Ć�<���<Ն�<Ɇ�<܆�<���<ӆ�<��<؆�<��<ӆ�<���<܆�<Ɇ�<Ն�<���<Ć�<چ�<���<���<`   `   ���<ӆ�<ۆ�<���<ˆ�<��<��<���<
��<ʆ�<ц�<��<Ԇ�<��<ц�<ʆ�<
��<���<��<��<ˆ�<���<ۆ�<ӆ�<`   `   ؆�<��<���<���<��<��<��<Ȇ�<ӆ�<Ԇ�<���<���<���<���<���<Ԇ�<ӆ�<Ȇ�<��<��<��<���<���<��<`   `   +��<҆�<���<ކ�<���<ǆ�<��<ކ�<͆�<܆�<��<��<؆�<��<��<܆�<͆�<ކ�<��<ǆ�<���<ކ�<���<҆�<`   `   ن�<��<ن�<ӆ�<ˆ�<؆�<���<ʆ�<ǆ�<Ć�<���<���<���<���<���<Ć�<ǆ�<ʆ�<���<؆�<ˆ�<ӆ�<ن�<��<`   `   ���<3��<8��<���<��<Æ�<���<���<Ć�<܆�<���<���<��<���<���<܆�<Ć�<���<���<Æ�<��<���<8��<3��<`   `   ���<@��<��<���<=��<]��<'��<"��<��<��<	��<��<U��<��<	��<��<��<"��<'��<]��<=��<���<��<@��<`   `   L��<.��<a��<N��<$��<G��</��<7��<.��<��<��<2��<\��<2��<��<��<.��<7��</��<G��<$��<N��<a��<.��<`   `   ��<��<e��<C��<!��<G��<��<1��<(��<C��<d��<`��<L��<`��<d��<C��<(��<1��<��<G��<!��<C��<e��<��<`   `   K��<��<��<��<t��<q��<��<H��<'��<��<,��<.��<��<.��<,��<��<'��<H��<��<q��<t��<��<��<��<`   `   ���<I��<H��<9��<k��<*��< ��<^��<%��<	��<��<(��<��<(��<��<	��<%��<^��< ��<*��<k��<9��<H��<I��<`   `   +��<,��<a��<B��<1��< ��<��<I��<��<A��<N��<?��<,��<?��<N��<A��<��<I��<��< ��<1��<B��<a��<,��<`   `   0��<=��<G��<��<:��<3��<?��<1��<��<f��<D��</��<<��</��<D��<f��<��<1��<?��<3��<:��<��<G��<=��<`   `   $��<7��<<��<��<+��</��<,��<��<"��<\��<��<,��<W��<,��<��<\��<"��<��<,��</��<+��<��<<��<7��<`   `   ��<��<P��<%��<��<2��<6��<��<��<;��<��<;��<[��<;��<��<;��<��<��<6��<2��<��<%��<P��<��<`   `   '��<4��<g��<2��<,��<,��<;��<_��<0��<-��<:��<N��<D��<N��<:��<-��<0��<_��<;��<,��<,��<2��<g��<4��<`   `   ��<'��<P��<8��<X��<��<��<c��<��<��<@��<7��<���<7��<@��<��<��<c��<��<��<X��<8��<P��<'��<`   `   7��<C��<;��<<��<���<2��<*��<Y��<��<���<-��<O��<%��<O��<-��<���<��<Y��<*��<2��<���<<��<;��<C��<`   `   N��<[��<2��<)��<[��<H��<n��<`��<c��<F��<��<b��<a��<b��<��<F��<c��<`��<n��<H��<[��<)��<2��<[��<`   `   ��<;��<0��<,��<��<��<K��<��<B��<Q��<���<��<��<��<���<Q��<B��<��<K��<��<��<,��<0��<;��<`   `   D��<0��< ��<<��<,��<K��<i��<���<��<3��<��<8��<4��<8��<��<3��<��<���<i��<K��<,��<<��< ��<0��<`   `   i��<#��<��<&��<(��<[��<w��<3��<.��<0��<.��<g��<w��<g��<.��<0��<.��<3��<w��<[��<(��<&��<��<#��<`   `   c��<?��<!��<"��<*��<(��<C��<7��<��<7��<1��<��<��<��<1��<7��<��<7��<C��<(��<*��<"��<!��<?��<`   `   >��<N��<4��<.��<^��<9��<`��<]��<��<6��<<��<-��<5��<-��<<��<6��<��<]��<`��<9��<^��<.��<4��<N��<`   `   
��<%��<0��<:��<L��<4��<X��<R��<��<)��<5��<f��<���<f��<5��<)��<��<R��<X��<4��<L��<:��<0��<%��<`   `   )��<#��<C��<H��<��<&��<+��<-��<D��<I��<M��<:��<+��<:��<M��<I��<D��<-��<+��<&��<��<H��<C��<#��<`   `   K��<*��<-��<7��<+��<3��<��<,��<4��<:��<;��<!��<:��<!��<;��<:��<4��<,��<��<3��<+��<7��<-��<*��<`   `   )��<-��<-��<2��<]��<C��<��<4��<��<<��<��<��<���<��<��<<��<��<4��<��<C��<]��<2��<-��<-��<`   `   ��<M��<u��<H��<R��<R��<C��<J��<:��<���<1��<��<H��<��<1��<���<:��<J��<C��<R��<R��<H��<u��<M��<`   `   H��<P��<r��<A��<��<-��<7��<O��<@��<7��<��<��<M��<��<��<7��<@��<O��<7��<-��<��<A��<r��<P��<`   `   U��<��<	��<��<��<"��<'��<]��<=��<���<��<@��<���<@��<��<���<=��<]��<'��<"��<��<��<	��<��<`   `   \��<2��<��<��<.��<7��</��<G��<$��<N��<a��<.��<L��<.��<a��<N��<$��<G��</��<7��<.��<��<��<2��<`   `   L��<`��<d��<C��<(��<1��<��<G��<!��<C��<e��<��<��<��<e��<C��<!��<G��<��<1��<(��<C��<d��<`��<`   `   ��<.��<,��<��<'��<H��<��<q��<t��<��<��<��<K��<��<��<��<t��<q��<��<H��<'��<��<,��<.��<`   `   ��<(��<��<	��<%��<^��< ��<*��<k��<9��<H��<I��<���<I��<H��<9��<k��<*��< ��<^��<%��<	��<��<(��<`   `   ,��<?��<N��<A��<��<I��<��< ��<1��<B��<a��<,��<+��<,��<a��<B��<1��< ��<��<I��<��<A��<N��<?��<`   `   <��</��<D��<f��<��<1��<?��<3��<:��<��<G��<=��<0��<=��<G��<��<:��<3��<?��<1��<��<f��<D��</��<`   `   W��<,��<��<\��<"��<��<,��</��<+��<��<<��<7��<$��<7��<<��<��<+��</��<,��<��<"��<\��<��<,��<`   `   [��<;��<��<;��<��<��<6��<2��<��<%��<P��<��<��<��<P��<%��<��<2��<6��<��<��<;��<��<;��<`   `   D��<N��<:��<-��<0��<_��<;��<,��<,��<2��<g��<4��<'��<4��<g��<2��<,��<,��<;��<_��<0��<-��<:��<N��<`   `   ���<7��<@��<��<��<c��<��<��<X��<8��<P��<'��<��<'��<P��<8��<X��<��<��<c��<��<��<@��<7��<`   `   %��<O��<-��<���<��<Y��<*��<2��<���<<��<;��<C��<7��<C��<;��<<��<���<2��<*��<Y��<��<���<-��<O��<`   `   a��<b��<��<F��<c��<`��<n��<H��<[��<)��<2��<[��<N��<[��<2��<)��<[��<H��<n��<`��<c��<F��<��<b��<`   `   ��<��<���<Q��<B��<��<K��<��<��<,��<0��<;��<��<;��<0��<,��<��<��<K��<��<B��<Q��<���<��<`   `   4��<8��<��<3��<��<���<i��<K��<,��<<��< ��<0��<D��<0��< ��<<��<,��<K��<i��<���<��<3��<��<8��<`   `   w��<g��<.��<0��<.��<3��<w��<[��<(��<&��<��<#��<i��<#��<��<&��<(��<[��<w��<3��<.��<0��<.��<g��<`   `   ��<��<1��<7��<��<7��<C��<(��<*��<"��<!��<?��<c��<?��<!��<"��<*��<(��<C��<7��<��<7��<1��<��<`   `   5��<-��<<��<6��<��<]��<`��<9��<^��<.��<4��<N��<>��<N��<4��<.��<^��<9��<`��<]��<��<6��<<��<-��<`   `   ���<f��<5��<)��<��<R��<X��<4��<L��<:��<0��<%��<
��<%��<0��<:��<L��<4��<X��<R��<��<)��<5��<f��<`   `   +��<:��<M��<I��<D��<-��<+��<&��<��<H��<C��<#��<)��<#��<C��<H��<��<&��<+��<-��<D��<I��<M��<:��<`   `   :��<!��<;��<:��<4��<,��<��<3��<+��<7��<-��<*��<K��<*��<-��<7��<+��<3��<��<,��<4��<:��<;��<!��<`   `   ���<��<��<<��<��<4��<��<C��<]��<2��<-��<-��<)��<-��<-��<2��<]��<C��<��<4��<��<<��<��<��<`   `   H��<��<1��<���<:��<J��<C��<R��<R��<H��<u��<M��<��<M��<u��<H��<R��<R��<C��<J��<:��<���<1��<��<`   `   M��<��<��<7��<@��<O��<7��<-��<��<A��<r��<P��<H��<P��<r��<A��<��<-��<7��<O��<@��<7��<��<��<`   `   h��<���<͉�<���<���<|��<���<z��<���<���<���<���<���<���<���<���<���<z��<���<|��<���<���<͉�<���<`   `   j��<���<���<���<���<���<���<���<ǉ�<���<���<���<U��<���<���<���<ǉ�<���<���<���<���<���<���<���<`   `   ���<ډ�<c��<e��<���<���<Ɖ�<���<ɉ�<���<���<���<{��<���<���<���<ɉ�<���<Ɖ�<���<���<e��<c��<ډ�<`   `   ���<��<���<���<���<Z��<���<���<���<���<���<���<��<���<���<���<���<���<���<Z��<���<���<���<��<`   `   r��<��<���<���<r��<���<͉�<���<���<���<���<t��<���<t��<���<���<���<���<͉�<���<r��<���<���<��<`   `   ���<Y��<x��<���<���<ɉ�<���<���<���<���<���<���<���<���<���<���<���<���<���<ɉ�<���<���<x��<Y��<`   `   ��<���<���<���<���<ȉ�<p��<���<���<m��<h��<ˉ�<���<ˉ�<h��<m��<���<���<p��<ȉ�<���<���<���<���<`   `   �<f��<͉�<���<���<É�<���<ɉ�<Չ�<���<t��<���<a��<���<t��<���<Չ�<ɉ�<���<É�<���<���<͉�<f��<`   `   ��<g��<���<ʉ�<���<���<���<���<���<���<���<���<��<���<���<���<���<���<���<���<���<ʉ�<���<g��<`   `   ��<���<z��<���<���<���<���<���<~��<���<���<̉�<v��<̉�<���<���<~��<���<���<���<���<���<z��<���<`   `   ���<���<}��<p��<���<���<���<���<��<���<���<���<���<���<���<���<��<���<���<���<���<p��<}��<���<`   `   n��<���<���<���<���<���<���<Y��<މ�<ĉ�<���<���<E��<���<���<ĉ�<މ�<Y��<���<���<���<���<���<���<`   `   ���<���<z��<���<���<t��<���<]��<���<���<���<���<���<���<���<���<���<]��<���<t��<���<���<z��<���<`   `   ���<���<z��<���<���<j��<���<���<���<���<ȉ�<���<���<���<ȉ�<���<���<���<���<j��<���<���<z��<���<`   `   ���<���<���<݉�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<݉�<���<���<`   `   ���<���<Ή�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<Ή�<���<`   `   ���<���<���<���<���<���<}��<���<���<���<���<���<���<���<���<���<���<���<}��<���<���<���<���<���<`   `   ���<���<���<���<���<���<y��<���<���<���<���<���<{��<���<���<���<���<���<y��<���<���<���<���<���<`   `   ɉ�<���<���<���<���<���<l��<���<É�<���<���<y��<k��<y��<���<���<É�<���<l��<���<���<���<���<���<`   `   Չ�<���<���<���<n��<Ɖ�<���<t��<���<���<���<���<���<���<���<���<���<t��<���<Ɖ�<n��<���<���<���<`   `   ω�<���<���<���<���<��<���<���<���<a��<���<���<���<���<���<a��<���<���<���<��<���<���<���<���<`   `   ���<���<���<���<���<p��<m��<݉�<���<p��<��<���<T��<���<��<p��<���<݉�<m��<p��<���<���<���<���<`   `   y��<���<���<t��<���<���<w��<���<}��<y��<Ӊ�<���<���<���<Ӊ�<y��<}��<���<w��<���<���<t��<���<���<`   `   ���<���<���<���<���<߉�<ω�<s��<d��<���<���<���<���<���<���<���<d��<s��<ω�<߉�<���<���<���<���<`   `   ���<���<���<���<���<z��<���<|��<���<���<͉�<���<h��<���<͉�<���<���<|��<���<z��<���<���<���<���<`   `   U��<���<���<���<ǉ�<���<���<���<���<���<���<���<j��<���<���<���<���<���<���<���<ǉ�<���<���<���<`   `   {��<���<���<���<ɉ�<���<Ɖ�<���<���<e��<c��<ډ�<���<ډ�<c��<e��<���<���<Ɖ�<���<ɉ�<���<���<���<`   `   ��<���<���<���<���<���<���<Z��<���<���<���<��<���<��<���<���<���<Z��<���<���<���<���<���<���<`   `   ���<t��<���<���<���<���<͉�<���<r��<���<���<��<r��<��<���<���<r��<���<͉�<���<���<���<���<t��<`   `   ���<���<���<���<���<���<���<ɉ�<���<���<x��<Y��<���<Y��<x��<���<���<ɉ�<���<���<���<���<���<���<`   `   ���<ˉ�<h��<m��<���<���<p��<ȉ�<���<���<���<���<��<���<���<���<���<ȉ�<p��<���<���<m��<h��<ˉ�<`   `   a��<���<t��<���<Չ�<ɉ�<���<É�<���<���<͉�<f��<�<f��<͉�<���<���<É�<���<ɉ�<Չ�<���<t��<���<`   `   ��<���<���<���<���<���<���<���<���<ʉ�<���<g��<��<g��<���<ʉ�<���<���<���<���<���<���<���<���<`   `   v��<̉�<���<���<~��<���<���<���<���<���<z��<���<��<���<z��<���<���<���<���<���<~��<���<���<̉�<`   `   ���<���<���<���<��<���<���<���<���<p��<}��<���<���<���<}��<p��<���<���<���<���<��<���<���<���<`   `   E��<���<���<ĉ�<މ�<Y��<���<���<���<���<���<���<n��<���<���<���<���<���<���<Y��<މ�<ĉ�<���<���<`   `   ���<���<���<���<���<]��<���<t��<���<���<z��<���<���<���<z��<���<���<t��<���<]��<���<���<���<���<`   `   ���<���<ȉ�<���<���<���<���<j��<���<���<z��<���<���<���<z��<���<���<j��<���<���<���<���<ȉ�<���<`   `   ���<���<���<���<���<���<���<���<���<݉�<���<���<���<���<���<݉�<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<Ή�<���<���<���<Ή�<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<���<���<}��<���<���<���<���<���<���<���<���<���<���<���<}��<���<���<���<���<���<`   `   {��<���<���<���<���<���<y��<���<���<���<���<���<���<���<���<���<���<���<y��<���<���<���<���<���<`   `   k��<y��<���<���<É�<���<l��<���<���<���<���<���<ɉ�<���<���<���<���<���<l��<���<É�<���<���<y��<`   `   ���<���<���<���<���<t��<���<Ɖ�<n��<���<���<���<Չ�<���<���<���<n��<Ɖ�<���<t��<���<���<���<���<`   `   ���<���<���<a��<���<���<���<��<���<���<���<���<ω�<���<���<���<���<��<���<���<���<a��<���<���<`   `   T��<���<��<p��<���<݉�<m��<p��<���<���<���<���<���<���<���<���<���<p��<m��<݉�<���<p��<��<���<`   `   ���<���<Ӊ�<y��<}��<���<w��<���<���<t��<���<���<y��<���<���<t��<���<���<w��<���<}��<y��<Ӊ�<���<`   `   ���<���<���<���<d��<s��<ω�<߉�<���<���<���<���<���<���<���<���<���<߉�<ω�<s��<d��<���<���<���<`   `   ��<��< ��<��<��<��<��<��<��<:��<1��< ��<��< ��<1��<:��<��<��<��<��<��<��< ��<��<`   `   
��<B��<��<��<��<��<��<��<
��<��<8��<,��<��<,��<8��<��<
��<��<��<��<��<��<��<B��<`   `   ��<2��<Պ�<L��<Z��<��<+��<���<��<��<���<���< ��<���<���<��<��<���<+��<��<Z��<L��<Պ�<2��<`   `   ���< ��<���<S��<��<��<"��<��<)��<��<��<��<*��<��<��<��<)��<��<"��<��<��<S��<���< ��<`   `   ���<��< ��<��<���<>��<#��<��<'��<���<��<��<3��<��<��<���<'��<��<#��<>��<���<��< ��<��<`   `   T��<F��<$��<,��<%��<��<���<��<-��<���<��<��<��<��<��<���<-��<��<���<��<%��<,��<$��<F��<`   `   
��< ��<��<��<��<Ԋ�<��<��<��<��<��<��<���<��<��<��<��<��<��<Ԋ�<��<��<��< ��<`   `   ��<���<��<��<��<��<!��<��<��<��<!��<L��<��<L��<!��<��<��<��<!��<��<��<��<��<���<`   `   "��<��<��<��<'��<��<��<��<���<#��<��<5��<U��<5��<��<#��<���<��<��<��<'��<��<��<��<`   `   ��<��<��<��<)��<��<��<��<��<��<ˊ�<��<6��<��<ˊ�<��<��<��<��<��<)��<��<��<��<`   `   ��<0��<8��<:��<��<-��<C��<��<���<��<��<��<i��<��<��<��<���<��<C��<-��<��<:��<8��<0��<`   `    ��<��<��<B��<ي�<���<8��<���<��<��<!��<��<G��<��<!��<��<��<���<8��<���<ي�<B��<��<��<`   `   ݊�<��<��<<��<��<&��<��<��<���<��<��<ي�<��<ي�<��<��<���<��<��<&��<��<<��<��<��<`   `   (��<,��<-��<���<+��<h��< ��<D��<��<���<��<���<L��<���<��<���<��<D��< ��<h��<+��<���<-��<,��<`   `   8��<*��<��<���< ��</��<Ҋ�<<��<��<���<7��<��<7��<��<7��<���<��<<��<Ҋ�</��< ��<���<��<*��<`   `   ��<��<���<��<%��<#��<���<'��<��<���<��<���<��<���<��<���<��<'��<���<#��<%��<��<���<��<`   `   ���<��<��<$��<,��<A��<F��< ��<(��< ��<��<��<-��<��<��< ��<(��< ��<F��<A��<,��<$��<��<��<`   `   ��<��<��<���<��</��<,��<���<��<��<��<8��<B��<8��<��<��<��<���<,��</��<��<���<��<��<`   `    ��<*��<��<��<���<1��<+��<&��<��<��<+��<��<��<��<+��<��<��<&��<+��<1��<���<��<��<*��<`   `   ��<��<��<��<��<��<��< ��<���<$��<��<#��<Y��<#��<��<$��<���< ��<��<��<��<��<��<��<`   `   ���<��< ��<��<��<���<��<��<���<9��<���<��<K��<��<���<9��<���<��<��<���<��<��< ��<��<`   `   ��</��<8��<E��<��<#��<@��<��<9��<0��<���<���<ϊ�<���<���<0��<9��<��<@��<#��<��<E��<8��</��<`   `   A��<"��<��<9��<��<��<��<��<C��<ي�<͊�<"��<$��<"��<͊�<ي�<C��<��<��<��<��<9��<��<"��<`   `   ��<��<��<!��<��<���<��<3��<B��<��<��< ��<6��< ��<��<��<B��<3��<��<���<��<!��<��<��<`   `   ��< ��<1��<:��<��<��<��<��<��<��< ��<��<��<��< ��<��<��<��<��<��<��<:��<1��< ��<`   `   ��<,��<8��<��<
��<��<��<��<��<��<��<B��<
��<B��<��<��<��<��<��<��<
��<��<8��<,��<`   `    ��<���<���<��<��<���<+��<��<Z��<L��<Պ�<2��<��<2��<Պ�<L��<Z��<��<+��<���<��<��<���<���<`   `   *��<��<��<��<)��<��<"��<��<��<S��<���< ��<���< ��<���<S��<��<��<"��<��<)��<��<��<��<`   `   3��<��<��<���<'��<��<#��<>��<���<��< ��<��<���<��< ��<��<���<>��<#��<��<'��<���<��<��<`   `   ��<��<��<���<-��<��<���<��<%��<,��<$��<F��<T��<F��<$��<,��<%��<��<���<��<-��<���<��<��<`   `   ���<��<��<��<��<��<��<Ԋ�<��<��<��< ��<
��< ��<��<��<��<Ԋ�<��<��<��<��<��<��<`   `   ��<L��<!��<��<��<��<!��<��<��<��<��<���<��<���<��<��<��<��<!��<��<��<��<!��<L��<`   `   U��<5��<��<#��<���<��<��<��<'��<��<��<��<"��<��<��<��<'��<��<��<��<���<#��<��<5��<`   `   6��<��<ˊ�<��<��<��<��<��<)��<��<��<��<��<��<��<��<)��<��<��<��<��<��<ˊ�<��<`   `   i��<��<��<��<���<��<C��<-��<��<:��<8��<0��<��<0��<8��<:��<��<-��<C��<��<���<��<��<��<`   `   G��<��<!��<��<��<���<8��<���<ي�<B��<��<��< ��<��<��<B��<ي�<���<8��<���<��<��<!��<��<`   `   ��<ي�<��<��<���<��<��<&��<��<<��<��<��<݊�<��<��<<��<��<&��<��<��<���<��<��<ي�<`   `   L��<���<��<���<��<D��< ��<h��<+��<���<-��<,��<(��<,��<-��<���<+��<h��< ��<D��<��<���<��<���<`   `   7��<��<7��<���<��<<��<Ҋ�</��< ��<���<��<*��<8��<*��<��<���< ��</��<Ҋ�<<��<��<���<7��<��<`   `   ��<���<��<���<��<'��<���<#��<%��<��<���<��<��<��<���<��<%��<#��<���<'��<��<���<��<���<`   `   -��<��<��< ��<(��< ��<F��<A��<,��<$��<��<��<���<��<��<$��<,��<A��<F��< ��<(��< ��<��<��<`   `   B��<8��<��<��<��<���<,��</��<��<���<��<��<��<��<��<���<��</��<,��<���<��<��<��<8��<`   `   ��<��<+��<��<��<&��<+��<1��<���<��<��<*��< ��<*��<��<��<���<1��<+��<&��<��<��<+��<��<`   `   Y��<#��<��<$��<���< ��<��<��<��<��<��<��<��<��<��<��<��<��<��< ��<���<$��<��<#��<`   `   K��<��<���<9��<���<��<��<���<��<��< ��<��<���<��< ��<��<��<���<��<��<���<9��<���<��<`   `   ϊ�<���<���<0��<9��<��<@��<#��<��<E��<8��</��<��</��<8��<E��<��<#��<@��<��<9��<0��<���<���<`   `   $��<"��<͊�<ي�<C��<��<��<��<��<9��<��<"��<A��<"��<��<9��<��<��<��<��<C��<ي�<͊�<"��<`   `   6��< ��<��<��<B��<3��<��<���<��<!��<��<��<��<��<��<!��<��<���<��<3��<B��<��<��< ��<`   `   �<v��<���<u��<v��<���<���<��<���<d��<o��<n��<��<n��<o��<d��<���<��<���<���<v��<u��<���<v��<`   `   ���<���<���<���<z��<���<���<ǌ�<���<���<v��<y��<ٌ�<y��<v��<���<���<ǌ�<���<���<z��<���<���<���<`   `   {��<���<���<���<a��<���<x��<���<���<���<���<���<݌�<���<���<���<���<���<x��<���<a��<���<���<���<`   `   ���<���<|��<r��<G��<���<���<���<ʌ�<���<݌�<���<_��<���<݌�<���<ʌ�<���<���<���<G��<r��<|��<���<`   `   ���<���<y��<���<���<���<g��<���<���<F��<���<���<r��<���<���<F��<���<���<g��<���<���<���<y��<���<`   `   O��<���<���<���<���<w��<���<���<���<y��<���<���<ڌ�<���<���<y��<���<���<���<w��<���<���<���<���<`   `   :��<���<v��<���<���<���<��<���<���<��<���<���<���<���<���<��<���<���<��<���<���<���<v��<���<`   `   ���<ʌ�<���<���<ʌ�<���<���<b��<g��<���<g��<_��<|��<_��<g��<���<g��<b��<���<���<ʌ�<���<���<ʌ�<`   `   ���<ˌ�<���<���<���<���<x��<���<���<���<���<���<���<���<���<���<���<���<x��<���<���<���<���<ˌ�<`   `   -��<���<���<~��<z��<���<���<ߌ�<���<���<��<r��<p��<r��<��<���<���<ߌ�<���<���<z��<~��<���<���<`   `   ���<���<n��<���<���<���<\��<���<i��<e��<��<o��<\��<o��<��<e��<i��<���<\��<���<���<���<n��<���<`   `   ��<���<C��<���<���<���<t��<��<���<e��<Ō�<���<���<���<Ō�<e��<���<��<t��<���<���<���<C��<���<`   `   ���<���<���<���<���<���<p��<Ō�<���<���<���<���<���<���<���<���<���<Ō�<p��<���<���<���<���<���<`   `   ���<���<Ȍ�<���<n��<���<r��<d��<���<Č�<���<f��<���<f��<���<Č�<���<d��<r��<���<n��<���<Ȍ�<���<`   `   u��<]��<���<ƌ�<��<���<���<w��<���<���<u��<���<���<���<u��<���<���<w��<���<���<��<ƌ�<���<]��<`   `   ���<���<���<̌�<���<l��<���<���<o��<���<���<���<���<���<���<���<o��<���<���<l��<���<̌�<���<���<`   `   ���<���<r��<���<���<V��<���<��<���<���<���<���<_��<���<���<���<���<��<���<V��<���<���<r��<���<`   `   ���<���<���<���<}��<c��<u��<i��<���<�<���<y��<���<y��<���<�<���<i��<u��<c��<}��<���<���<���<`   `   q��<}��<���<̌�<ʌ�<���<���<���<���<���<���<���<~��<���<���<���<���<���<���<���<ʌ�<̌�<���<}��<`   `   ���<���<���<���<��<k��<~��<܌�<���<���<���<q��<]��<q��<���<���<���<܌�<~��<k��<��<���<���<���<`   `   ���<ǌ�<~��<i��<���<=��<w��<���<���<���<w��<���<���<���<w��<���<���<���<w��<=��<���<i��<~��<ǌ�<`   `   q��<z��<^��<g��<���<���<֌�<e��<m��<���<���<���<���<���<���<���<m��<e��<֌�<���<���<g��<^��<z��<`   `   ���<���<���<���<���<���<���<g��<���<ʌ�<Ȍ�<���<���<���<Ȍ�<ʌ�<���<g��<���<���<���<���<���<���<`   `   ���<���<���<���<���<���<k��<���<���<���<���<i��<���<i��<���<���<���<���<k��<���<���<���<���<���<`   `   ��<n��<o��<d��<���<��<���<���<v��<u��<���<v��<�<v��<���<u��<v��<���<���<��<���<d��<o��<n��<`   `   ٌ�<y��<v��<���<���<ǌ�<���<���<z��<���<���<���<���<���<���<���<z��<���<���<ǌ�<���<���<v��<y��<`   `   ݌�<���<���<���<���<���<x��<���<a��<���<���<���<{��<���<���<���<a��<���<x��<���<���<���<���<���<`   `   _��<���<݌�<���<ʌ�<���<���<���<G��<r��<|��<���<���<���<|��<r��<G��<���<���<���<ʌ�<���<݌�<���<`   `   r��<���<���<F��<���<���<g��<���<���<���<y��<���<���<���<y��<���<���<���<g��<���<���<F��<���<���<`   `   ڌ�<���<���<y��<���<���<���<w��<���<���<���<���<O��<���<���<���<���<w��<���<���<���<y��<���<���<`   `   ���<���<���<��<���<���<��<���<���<���<v��<���<:��<���<v��<���<���<���<��<���<���<��<���<���<`   `   |��<_��<g��<���<g��<b��<���<���<ʌ�<���<���<ʌ�<���<ʌ�<���<���<ʌ�<���<���<b��<g��<���<g��<_��<`   `   ���<���<���<���<���<���<x��<���<���<���<���<ˌ�<���<ˌ�<���<���<���<���<x��<���<���<���<���<���<`   `   p��<r��<��<���<���<ߌ�<���<���<z��<~��<���<���<-��<���<���<~��<z��<���<���<ߌ�<���<���<��<r��<`   `   \��<o��<��<e��<i��<���<\��<���<���<���<n��<���<���<���<n��<���<���<���<\��<���<i��<e��<��<o��<`   `   ���<���<Ō�<e��<���<��<t��<���<���<���<C��<���<��<���<C��<���<���<���<t��<��<���<e��<Ō�<���<`   `   ���<���<���<���<���<Ō�<p��<���<���<���<���<���<���<���<���<���<���<���<p��<Ō�<���<���<���<���<`   `   ���<f��<���<Č�<���<d��<r��<���<n��<���<Ȍ�<���<���<���<Ȍ�<���<n��<���<r��<d��<���<Č�<���<f��<`   `   ���<���<u��<���<���<w��<���<���<��<ƌ�<���<]��<u��<]��<���<ƌ�<��<���<���<w��<���<���<u��<���<`   `   ���<���<���<���<o��<���<���<l��<���<̌�<���<���<���<���<���<̌�<���<l��<���<���<o��<���<���<���<`   `   _��<���<���<���<���<��<���<V��<���<���<r��<���<���<���<r��<���<���<V��<���<��<���<���<���<���<`   `   ���<y��<���<�<���<i��<u��<c��<}��<���<���<���<���<���<���<���<}��<c��<u��<i��<���<�<���<y��<`   `   ~��<���<���<���<���<���<���<���<ʌ�<̌�<���<}��<q��<}��<���<̌�<ʌ�<���<���<���<���<���<���<���<`   `   ]��<q��<���<���<���<܌�<~��<k��<��<���<���<���<���<���<���<���<��<k��<~��<܌�<���<���<���<q��<`   `   ���<���<w��<���<���<���<w��<=��<���<i��<~��<ǌ�<���<ǌ�<~��<i��<���<=��<w��<���<���<���<w��<���<`   `   ���<���<���<���<m��<e��<֌�<���<���<g��<^��<z��<q��<z��<^��<g��<���<���<֌�<e��<m��<���<���<���<`   `   ���<���<Ȍ�<ʌ�<���<g��<���<���<���<���<���<���<���<���<���<���<���<���<���<g��<���<ʌ�<Ȍ�<���<`   `   ���<i��<���<���<���<���<k��<���<���<���<���<���<���<���<���<���<���<���<k��<���<���<���<���<i��<`   `   ��<��<��<)��<+��<��<��<��<��<8��<C��<J��<��<J��<C��<8��<��<��<��<��<+��<)��<��<��<`   `   4��<���<$��<,��<h��<A��<��<��<��<o��<=��<��<	��<��<=��<o��<��<��<��<A��<h��<,��<$��<���<`   `   0��<��<*��<���<(��<Q��<!��<��<��<0��<��<��<(��<��<��<0��<��<��<!��<Q��<(��<���<*��<��<`   `   V��<#��<7��<1��<,��<?��<)��<*��<��<��<��<#��<X��<#��<��<��<��<*��<)��<?��<,��<1��<7��<#��<`   `   ��<��<0��<c��<M��<"��<#��<5��<%��<a��<>��<��<4��<��<>��<a��<%��<5��<#��<"��<M��<c��<0��<��<`   `   ��<(��<��<
��<
��<��<'��<��<��<?��<��<��<5��<��<��<?��<��<��<'��<��<
��<
��<��<(��<`   `   m��<^��<"��<��<��<*��<��<��<'��<���<��<2��<V��<2��<��<���<'��<��<��<*��<��<��<"��<^��<`   `   .��<��<���<J��<��<��<��<��<p��<��<>��<H��<%��<H��<>��<��<p��<��<��<��<��<J��<���<��<`   `   &��<���<��<C��<��<;��<+��<��<+��<��<9��<2��<��<2��<9��<��<+��<��<+��<;��<��<C��<��<���<`   `   w��<A��<��<I��<��<l��<Y��<��<��<��<2��<A��<X��<A��<2��<��<��<��<Y��<l��<��<I��<��<A��<`   `   '��</��<-��<4��<��<>��<��<��<E��<'��<��<(��<_��<(��<��<'��<E��<��<��<>��<��<4��<-��</��<`   `   ���<��<_��<"��<(��<W��<+��<��<D��<+��<��<���<&��<���<��<+��<D��<��<+��<W��<(��<"��<_��<��<`   `   ���<<��<T��<��<*��<"��<4��<���<��<��<��<H��<%��<H��<��<��<��<���<4��<"��<*��<��<T��<<��<`   `   T��<��<��<&��<-��<���<T��<(��<	��<��<*��<c��<���<c��<*��<��<	��<(��<T��<���<-��<&��<��<��<`   `   U��<!��<��<B��<B��<#��<d��<E��<l��<5��<��<7��<ލ�<7��<��<5��<l��<E��<d��<#��<B��<B��<��<!��<`   `   ��<Z��<O��<���< ��<��<��<��<G��<(��<��<D��<(��<D��<��<(��<G��<��<��<��< ��<���<O��<Z��<`   `   ύ�<&��<��<��<I��<L��</��<>��<��<���<��<,��<2��<,��<��<���<��<>��</��<L��<I��<��<��<&��<`   `   7��<0��<)��<.��<<��<U��<;��<I��<.��<��<��<%��<O��<%��<��<��<.��<I��<;��<U��<<��<.��<)��<0��<`   `   o��<%��<"��<��<č�<4��<��<���<%��<��<��<=��<p��<=��<��<��<%��<���<��<4��<č�<��<"��<%��<`   `   2��<���<"��<���<��<c��<8��<���<��<��<*��<;��<��<;��<*��<��<��<���<8��<c��<��<���<"��<���<`   `   N��<$��<i��<P��<<��<_��</��<?��<E��<��<9��<J��<���<J��<9��<��<E��<?��</��<_��<<��<P��<i��<$��<`   `   G��<��<E��<6��< ��<��<	��<a��<<��<���<��<B��<��<B��<��<���<<��<a��<	��<��< ��<6��<E��<��<`   `   ��<��<��<��<)��<���<��<\��<
��<��<��<��<��<��<��<��<
��<\��<��<���<)��<��<��<��<`   `   ��<@��<2��<(��<G��<$��<��<5��<��<��<3��<��<?��<��<3��<��<��<5��<��<$��<G��<(��<2��<@��<`   `   ��<J��<C��<8��<��<��<��<��<+��<)��<��<��<��<��<��<)��<+��<��<��<��<��<8��<C��<J��<`   `   	��<��<=��<o��<��<��<��<A��<h��<,��<$��<���<4��<���<$��<,��<h��<A��<��<��<��<o��<=��<��<`   `   (��<��<��<0��<��<��<!��<Q��<(��<���<*��<��<0��<��<*��<���<(��<Q��<!��<��<��<0��<��<��<`   `   X��<#��<��<��<��<*��<)��<?��<,��<1��<7��<#��<V��<#��<7��<1��<,��<?��<)��<*��<��<��<��<#��<`   `   4��<��<>��<a��<%��<5��<#��<"��<M��<c��<0��<��<��<��<0��<c��<M��<"��<#��<5��<%��<a��<>��<��<`   `   5��<��<��<?��<��<��<'��<��<
��<
��<��<(��<��<(��<��<
��<
��<��<'��<��<��<?��<��<��<`   `   V��<2��<��<���<'��<��<��<*��<��<��<"��<^��<m��<^��<"��<��<��<*��<��<��<'��<���<��<2��<`   `   %��<H��<>��<��<p��<��<��<��<��<J��<���<��<.��<��<���<J��<��<��<��<��<p��<��<>��<H��<`   `   ��<2��<9��<��<+��<��<+��<;��<��<C��<��<���<&��<���<��<C��<��<;��<+��<��<+��<��<9��<2��<`   `   X��<A��<2��<��<��<��<Y��<l��<��<I��<��<A��<w��<A��<��<I��<��<l��<Y��<��<��<��<2��<A��<`   `   _��<(��<��<'��<E��<��<��<>��<��<4��<-��</��<'��</��<-��<4��<��<>��<��<��<E��<'��<��<(��<`   `   &��<���<��<+��<D��<��<+��<W��<(��<"��<_��<��<���<��<_��<"��<(��<W��<+��<��<D��<+��<��<���<`   `   %��<H��<��<��<��<���<4��<"��<*��<��<T��<<��<���<<��<T��<��<*��<"��<4��<���<��<��<��<H��<`   `   ���<c��<*��<��<	��<(��<T��<���<-��<&��<��<��<T��<��<��<&��<-��<���<T��<(��<	��<��<*��<c��<`   `   ލ�<7��<��<5��<l��<E��<d��<#��<B��<B��<��<!��<U��<!��<��<B��<B��<#��<d��<E��<l��<5��<��<7��<`   `   (��<D��<��<(��<G��<��<��<��< ��<���<O��<Z��<��<Z��<O��<���< ��<��<��<��<G��<(��<��<D��<`   `   2��<,��<��<���<��<>��</��<L��<I��<��<��<&��<ύ�<&��<��<��<I��<L��</��<>��<��<���<��<,��<`   `   O��<%��<��<��<.��<I��<;��<U��<<��<.��<)��<0��<7��<0��<)��<.��<<��<U��<;��<I��<.��<��<��<%��<`   `   p��<=��<��<��<%��<���<��<4��<č�<��<"��<%��<o��<%��<"��<��<č�<4��<��<���<%��<��<��<=��<`   `   ��<;��<*��<��<��<���<8��<c��<��<���<"��<���<2��<���<"��<���<��<c��<8��<���<��<��<*��<;��<`   `   ���<J��<9��<��<E��<?��</��<_��<<��<P��<i��<$��<N��<$��<i��<P��<<��<_��</��<?��<E��<��<9��<J��<`   `   ��<B��<��<���<<��<a��<	��<��< ��<6��<E��<��<G��<��<E��<6��< ��<��<	��<a��<<��<���<��<B��<`   `   ��<��<��<��<
��<\��<��<���<)��<��<��<��<��<��<��<��<)��<���<��<\��<
��<��<��<��<`   `   ?��<��<3��<��<��<5��<��<$��<G��<(��<2��<@��<��<@��<2��<(��<G��<$��<��<5��<��<��<3��<��<`   `   ���<ʏ�<���<���<͏�<���<��<���<���<���<���<��<ҏ�<��<���<���<���<���<��<���<͏�<���<���<ʏ�<`   `   ���<܏�<Տ�<���<���<���<��<Տ�<���<���<���<���<���<���<���<���<���<Տ�<��<���<���<���<Տ�<܏�<`   `   ���<�<ŏ�<���<ŏ�<���<ҏ�<���<��<ˏ�<���<��<t��<��<���<ˏ�<��<���<ҏ�<���<ŏ�<���<ŏ�<�<`   `   ď�<���<���<���<֏�<���<���<���<���<ď�<���<���<̏�<���<���<ď�<���<���<���<���<֏�<���<���<���<`   `   ��<�<�<���<���<���<ߏ�<ˏ�<���<��<���<ُ�<ڏ�<ُ�<���<��<���<ˏ�<ߏ�<���<���<���<�<�<`   `   ���<ˏ�<Ə�<���<���<֏�<ʏ�<؏�<ɏ�<Џ�<ҏ�<���<���<���<ҏ�<Џ�<ɏ�<؏�<ʏ�<֏�<���<���<Ə�<ˏ�<`   `   ���<���<ݏ�<��<��<���<���<Ǐ�<���<}��<ӏ�<Ǐ�<���<Ǐ�<ӏ�<}��<���<Ǐ�<���<���<��<��<ݏ�<���<`   `   ���<���<��<���<���<��<Џ�<��<ݏ�<���<���<ď�<���<ď�<���<���<ݏ�<��<Џ�<��<���<���<��<���<`   `   ���<��<��<���<���<Ǐ�<؏�<���<���<��<͏�<���<���<���<͏�<��<���<���<؏�<Ǐ�<���<���<��<��<`   `   ���<̏�<���<ߏ�<׏�<���<���<���<я�<׏�<���<���<���<���<���<׏�<я�<���<���<���<׏�<ߏ�<���<̏�<`   `   ���<���<���<Ǐ�<���<���<؏�<܏�<��<��<���<ڏ�<ď�<ڏ�<���<��<��<܏�<؏�<���<���<Ǐ�<���<���<`   `   ��<Ϗ�<Ώ�<���<���<���<���<���<���<��<Џ�<��<���<��<Џ�<��<���<���<���<���<���<���<Ώ�<Ϗ�<`   `   ���<ԏ�<ɏ�<���<��<���<֏�<ӏ�<ُ�<��<���<ŏ�<���<ŏ�<���<��<ُ�<ӏ�<֏�<���<��<���<ɏ�<ԏ�<`   `   ȏ�<ȏ�<���<���<���<���<���<��<ڏ�<���<���<��<���<��<���<���<ڏ�<��<���<���<���<���<���<ȏ�<`   `   ȏ�<ȏ�<ʏ�<���<ڏ�<Տ�<���<���<���<���<Ϗ�<��<���<��<Ϗ�<���<���<���<���<Տ�<ڏ�<���<ʏ�<ȏ�<`   `   ���<���<ݏ�<���<���<ڏ�<���<���<���<ُ�<���<���<ʏ�<���<���<ُ�<���<���<���<ڏ�<���<���<ݏ�<���<`   `   �<���<ݏ�<Џ�<ď�<ȏ�<���<��<���<ŏ�<��<���<͏�<���<��<ŏ�<���<��<���<ȏ�<ď�<Џ�<ݏ�<���<`   `   Ϗ�<Ǐ�<ȏ�<��<؏�<���<���<ݏ�<���<ď�<��<���<���<���<��<ď�<���<ݏ�<���<���<؏�<��<ȏ�<Ǐ�<`   `   ʏ�<ҏ�<׏�<���<ڏ�<���<���<Ώ�<��<ُ�<���<���<���<���<���<ُ�<��<Ώ�<���<���<ڏ�<���<׏�<ҏ�<`   `   ���<���<я�<��<���<���<ˏ�<���<ӏ�<ҏ�<���<���<̏�<���<���<ҏ�<ӏ�<���<ˏ�<���<���<��<я�<���<`   `   ���<���<���<���<���<Ώ�<���<���<���<ۏ�<̏�<���<���<���<̏�<ۏ�<���<���<���<Ώ�<���<���<���<���<`   `   ���<���<ڏ�<���<���<׏�<���<���<ʏ�<��<���<���<���<���<���<��<ʏ�<���<���<׏�<���<���<ڏ�<���<`   `   ���<ӏ�<͏�<���<̏�<��<Ə�<���<��<���<���<я�<���<я�<���<���<��<���<Ə�<��<̏�<���<͏�<ӏ�<`   `   ���<���<���<Ǐ�<ُ�<̏�<��<���<؏�<Џ�<���<ԏ�<���<ԏ�<���<Џ�<؏�<���<��<̏�<ُ�<Ǐ�<���<���<`   `   ҏ�<��<���<���<���<���<��<���<͏�<���<���<ʏ�<���<ʏ�<���<���<͏�<���<��<���<���<���<���<��<`   `   ���<���<���<���<���<Տ�<��<���<���<���<Տ�<܏�<���<܏�<Տ�<���<���<���<��<Տ�<���<���<���<���<`   `   t��<��<���<ˏ�<��<���<ҏ�<���<ŏ�<���<ŏ�<�<���<�<ŏ�<���<ŏ�<���<ҏ�<���<��<ˏ�<���<��<`   `   ̏�<���<���<ď�<���<���<���<���<֏�<���<���<���<ď�<���<���<���<֏�<���<���<���<���<ď�<���<���<`   `   ڏ�<ُ�<���<��<���<ˏ�<ߏ�<���<���<���<�<�<��<�<�<���<���<���<ߏ�<ˏ�<���<��<���<ُ�<`   `   ���<���<ҏ�<Џ�<ɏ�<؏�<ʏ�<֏�<���<���<Ə�<ˏ�<���<ˏ�<Ə�<���<���<֏�<ʏ�<؏�<ɏ�<Џ�<ҏ�<���<`   `   ���<Ǐ�<ӏ�<}��<���<Ǐ�<���<���<��<��<ݏ�<���<���<���<ݏ�<��<��<���<���<Ǐ�<���<}��<ӏ�<Ǐ�<`   `   ���<ď�<���<���<ݏ�<��<Џ�<��<���<���<��<���<���<���<��<���<���<��<Џ�<��<ݏ�<���<���<ď�<`   `   ���<���<͏�<��<���<���<؏�<Ǐ�<���<���<��<��<���<��<��<���<���<Ǐ�<؏�<���<���<��<͏�<���<`   `   ���<���<���<׏�<я�<���<���<���<׏�<ߏ�<���<̏�<���<̏�<���<ߏ�<׏�<���<���<���<я�<׏�<���<���<`   `   ď�<ڏ�<���<��<��<܏�<؏�<���<���<Ǐ�<���<���<���<���<���<Ǐ�<���<���<؏�<܏�<��<��<���<ڏ�<`   `   ���<��<Џ�<��<���<���<���<���<���<���<Ώ�<Ϗ�<��<Ϗ�<Ώ�<���<���<���<���<���<���<��<Џ�<��<`   `   ���<ŏ�<���<��<ُ�<ӏ�<֏�<���<��<���<ɏ�<ԏ�<���<ԏ�<ɏ�<���<��<���<֏�<ӏ�<ُ�<��<���<ŏ�<`   `   ���<��<���<���<ڏ�<��<���<���<���<���<���<ȏ�<ȏ�<ȏ�<���<���<���<���<���<��<ڏ�<���<���<��<`   `   ���<��<Ϗ�<���<���<���<���<Տ�<ڏ�<���<ʏ�<ȏ�<ȏ�<ȏ�<ʏ�<���<ڏ�<Տ�<���<���<���<���<Ϗ�<��<`   `   ʏ�<���<���<ُ�<���<���<���<ڏ�<���<���<ݏ�<���<���<���<ݏ�<���<���<ڏ�<���<���<���<ُ�<���<���<`   `   ͏�<���<��<ŏ�<���<��<���<ȏ�<ď�<Џ�<ݏ�<���<�<���<ݏ�<Џ�<ď�<ȏ�<���<��<���<ŏ�<��<���<`   `   ���<���<��<ď�<���<ݏ�<���<���<؏�<��<ȏ�<Ǐ�<Ϗ�<Ǐ�<ȏ�<��<؏�<���<���<ݏ�<���<ď�<��<���<`   `   ���<���<���<ُ�<��<Ώ�<���<���<ڏ�<���<׏�<ҏ�<ʏ�<ҏ�<׏�<���<ڏ�<���<���<Ώ�<��<ُ�<���<���<`   `   ̏�<���<���<ҏ�<ӏ�<���<ˏ�<���<���<��<я�<���<���<���<я�<��<���<���<ˏ�<���<ӏ�<ҏ�<���<���<`   `   ���<���<̏�<ۏ�<���<���<���<Ώ�<���<���<���<���<���<���<���<���<���<Ώ�<���<���<���<ۏ�<̏�<���<`   `   ���<���<���<��<ʏ�<���<���<׏�<���<���<ڏ�<���<���<���<ڏ�<���<���<׏�<���<���<ʏ�<��<���<���<`   `   ���<я�<���<���<��<���<Ə�<��<̏�<���<͏�<ӏ�<���<ӏ�<͏�<���<̏�<��<Ə�<���<��<���<���<я�<`   `   ���<ԏ�<���<Џ�<؏�<���<��<̏�<ُ�<Ǐ�<���<���<���<���<���<Ǐ�<ُ�<̏�<��<���<؏�<Џ�<���<ԏ�<`   `   2��<}��<^��<g��<���<t��<q��<k��<���<���<���<Z��<a��<Z��<���<���<���<k��<q��<t��<���<g��<^��<}��<`   `   x��<r��<l��<{��<g��<q��<t��<W��<b��<N��<S��<i��<f��<i��<S��<N��<b��<W��<t��<q��<g��<{��<l��<r��<`   `   y��<\��<v��<���<{��<{��<i��<H��<m��<{��<���<���<E��<���<���<{��<m��<H��<i��<{��<{��<���<v��<\��<`   `   W��<`��<p��<_��<���<���<t��<L��<���<���<v��<p��<	��<p��<v��<���<���<L��<t��<���<���<_��<p��<`��<`   `   q��<���<{��<I��<x��<z��<���<_��<N��<0��<0��<w��<3��<w��<0��<0��<N��<_��<���<z��<x��<I��<{��<���<`   `   T��<G��<q��<}��<}��<Z��<`��<x��<y��<k��<t��<���<���<���<t��<k��<y��<x��<`��<Z��<}��<}��<q��<G��<`   `   b��<6��<P��<e��<]��<H��<I��<i��<s��<���<n��<d��<���<d��<n��<���<s��<i��<I��<H��<]��<e��<P��<6��<`   `   ���<���<f��<J��<o��<j��<���<h��<#��<r��<-��<6��<���<6��<-��<r��<#��<h��<���<j��<o��<J��<f��<���<`   `   k��<���<p��<P��<���<^��<i��<g��<8��<���<a��<���<ߑ�<���<a��<���<8��<g��<i��<^��<���<P��<p��<���<`   `   ��<d��<h��<8��<���<[��<N��<���<u��<|��<���<���<t��<���<���<|��<u��<���<N��<[��<���<8��<h��<d��<`   `   ���<x��<���<`��<���<���<z��<���<5��<"��<���<x��<���<x��<���<"��<5��<���<z��<���<���<`��<���<x��<`   `   ߑ�<^��<U��<{��<���<w��<O��<`��<��<1��<���<���<S��<���<���<1��<��<`��<O��<w��<���<{��<U��<^��<`   `   x��<0��<N��<`��<m��<r��<I��<t��<���<���<L��<a��<���<a��<L��<���<���<t��<I��<r��<m��<`��<N��<0��<`   `   :��<{��<Ǒ�<k��<S��<���<d��<k��<s��<���<Q��<L��<���<L��<Q��<���<s��<k��<d��<���<S��<k��<Ǒ�<{��<`   `   b��<o��<���<~��<G��<x��<���<}��<8��<l��<���<^��<���<^��<���<l��<8��<}��<���<x��<G��<~��<���<o��<`   `   ���<-��<H��<Ñ�<r��<���<���<ő�<��<z��<j��<A��<���<A��<j��<z��<��<ő�<���<���<r��<Ñ�<H��<-��<`   `   ��<x��<o��<���<K��<g��<w��<t��<���<y��<N��<W��<���<W��<N��<y��<���<t��<w��<g��<K��<���<o��<x��<`   `   \��<s��<F��<+��<2��<g��<o��<5��<X��<\��<b��<���<���<���<b��<\��<X��<5��<o��<g��<2��<+��<F��<s��<`   `   ��<|��<B��<K��<���<|��<���<l��<b��<S��<l��<���<h��<���<l��<S��<b��<l��<���<|��<���<K��<B��<|��<`   `   ���<ߑ�<o��<p��<���<.��<v��<���<a��<U��<k��<���<���<���<k��<U��<a��<���<v��<.��<���<p��<o��<ߑ�<`   `   ���<���<K��<H��<q��<2��<���<���<L��<S��<d��<c��<���<c��<d��<S��<L��<���<���<2��<q��<H��<K��<���<`   `   N��<X��<n��<t��<���<���<���<���<?��<c��<k��<a��<���<a��<k��<c��<?��<���<���<���<���<t��<n��<X��<`   `   ]��<m��<���<e��<K��<b��<l��<H��<>��<_��<d��<x��<g��<x��<d��<_��<>��<H��<l��<b��<K��<e��<���<m��<`   `   g��<o��<���<���<Z��<B��<N��<B��<k��<T��<W��<���</��<���<W��<T��<k��<B��<N��<B��<Z��<���<���<o��<`   `   a��<Z��<���<���<���<k��<q��<t��<���<g��<^��<}��<2��<}��<^��<g��<���<t��<q��<k��<���<���<���<Z��<`   `   f��<i��<S��<N��<b��<W��<t��<q��<g��<{��<l��<r��<x��<r��<l��<{��<g��<q��<t��<W��<b��<N��<S��<i��<`   `   E��<���<���<{��<m��<H��<i��<{��<{��<���<v��<\��<y��<\��<v��<���<{��<{��<i��<H��<m��<{��<���<���<`   `   	��<p��<v��<���<���<L��<t��<���<���<_��<p��<`��<W��<`��<p��<_��<���<���<t��<L��<���<���<v��<p��<`   `   3��<w��<0��<0��<N��<_��<���<z��<x��<I��<{��<���<q��<���<{��<I��<x��<z��<���<_��<N��<0��<0��<w��<`   `   ���<���<t��<k��<y��<x��<`��<Z��<}��<}��<q��<G��<T��<G��<q��<}��<}��<Z��<`��<x��<y��<k��<t��<���<`   `   ���<d��<n��<���<s��<i��<I��<H��<]��<e��<P��<6��<b��<6��<P��<e��<]��<H��<I��<i��<s��<���<n��<d��<`   `   ���<6��<-��<r��<#��<h��<���<j��<o��<J��<f��<���<���<���<f��<J��<o��<j��<���<h��<#��<r��<-��<6��<`   `   ߑ�<���<a��<���<8��<g��<i��<^��<���<P��<p��<���<k��<���<p��<P��<���<^��<i��<g��<8��<���<a��<���<`   `   t��<���<���<|��<u��<���<N��<[��<���<8��<h��<d��<��<d��<h��<8��<���<[��<N��<���<u��<|��<���<���<`   `   ���<x��<���<"��<5��<���<z��<���<���<`��<���<x��<���<x��<���<`��<���<���<z��<���<5��<"��<���<x��<`   `   S��<���<���<1��<��<`��<O��<w��<���<{��<U��<^��<ߑ�<^��<U��<{��<���<w��<O��<`��<��<1��<���<���<`   `   ���<a��<L��<���<���<t��<I��<r��<m��<`��<N��<0��<x��<0��<N��<`��<m��<r��<I��<t��<���<���<L��<a��<`   `   ���<L��<Q��<���<s��<k��<d��<���<S��<k��<Ǒ�<{��<:��<{��<Ǒ�<k��<S��<���<d��<k��<s��<���<Q��<L��<`   `   ���<^��<���<l��<8��<}��<���<x��<G��<~��<���<o��<b��<o��<���<~��<G��<x��<���<}��<8��<l��<���<^��<`   `   ���<A��<j��<z��<��<ő�<���<���<r��<Ñ�<H��<-��<���<-��<H��<Ñ�<r��<���<���<ő�<��<z��<j��<A��<`   `   ���<W��<N��<y��<���<t��<w��<g��<K��<���<o��<x��<��<x��<o��<���<K��<g��<w��<t��<���<y��<N��<W��<`   `   ���<���<b��<\��<X��<5��<o��<g��<2��<+��<F��<s��<\��<s��<F��<+��<2��<g��<o��<5��<X��<\��<b��<���<`   `   h��<���<l��<S��<b��<l��<���<|��<���<K��<B��<|��<��<|��<B��<K��<���<|��<���<l��<b��<S��<l��<���<`   `   ���<���<k��<U��<a��<���<v��<.��<���<p��<o��<ߑ�<���<ߑ�<o��<p��<���<.��<v��<���<a��<U��<k��<���<`   `   ���<c��<d��<S��<L��<���<���<2��<q��<H��<K��<���<���<���<K��<H��<q��<2��<���<���<L��<S��<d��<c��<`   `   ���<a��<k��<c��<?��<���<���<���<���<t��<n��<X��<N��<X��<n��<t��<���<���<���<���<?��<c��<k��<a��<`   `   g��<x��<d��<_��<>��<H��<l��<b��<K��<e��<���<m��<]��<m��<���<e��<K��<b��<l��<H��<>��<_��<d��<x��<`   `   /��<���<W��<T��<k��<B��<N��<B��<Z��<���<���<o��<g��<o��<���<���<Z��<B��<N��<B��<k��<T��<W��<���<`   `   X��</��<��<7��<��<@��<	��<Q��<5��<��<W��<��<H��<��<W��<��<5��<Q��<	��<@��<��<7��<��</��<`   `   ?��<��<���<+��<��<H��<���<%��<��<��<D��<��<a��<��<D��<��<��<%��<���<H��<��<+��<���<��<`   `   F��<��<��<(��<��</��<��<0��<���<��<��< ��<���< ��<��<��<���<0��<��</��<��<(��<��<��<`   `   ��<*��<&��<��<���<	��<+��<Z��<4��<3��<&��< ��<t��< ��<&��<3��<4��<Z��<+��<	��<���<��<&��<*��<`   `   ��<��<��<$��</��<��<��<��<0��<9��<;��<7��<0��<7��<;��<9��<0��<��<��<��</��<$��<��<��<`   `   0��<7��<3��<9��<1��<,��<7��<��<��<&��<��<��<���<��<��<&��<��<��<7��<,��<1��<9��<3��<7��<`   `   W��<W��<>��<��<���<)��<O��< ��<%��<>��<��<��<#��<��<��<>��<%��< ��<O��<)��<���<��<>��<W��<`   `   ��<��<��<J��<:��<��<!��<'��<=��<5��<4��<8��<��<8��<4��<5��<=��<'��<!��<��<:��<J��<��<��<`   `   ��<ؒ�<��<a��<.��<��<)��<<��<N��<��<��<#��<���<#��<��<��<N��<<��<)��<��<.��<a��<��<ؒ�<`   `   |��<;��<E��<��<Ւ�<.��<@��<��<'��<��<
��<4��<���<4��<
��<��<'��<��<@��<.��<Ւ�<��<E��<;��<`   `   ��<%��<p��<��<��<M��<��<��<R��<`��<���<��<V��<��<���<`��<R��<��<��<M��<��<��<p��<%��<`   `   ��<��<j��<;��<���<��<���<V��<~��<h��<��<���<N��<���<��<h��<~��<V��<���<��<���<;��<j��<��<`   `   F��<2��<B��<?��<��<N��<D��<>��<��<��<F��<��<9��<��<F��<��<��<>��<D��<N��<��<?��<B��<2��<`   `   H��<A��<��</��<3��<`��<8��<��<��<��<C��<��<(��<��<C��<��<��<��<8��<`��<3��</��<��<A��<`   `   K��<X��<��<��<4��<��<���<6��<T��<$��<7��<��<��<��<7��<$��<T��<6��<���<��<4��<��<��<X��<`   `   ��<A��<���<��<1��<��<��<��<��<���<>��<3��<��<3��<>��<���<��<��<��<��<1��<��<���<A��<`   `   ے�<&��<G��<$��<@��<U��<��<ݒ�<%��<��<.��<<��<���<<��<.��<��<%��<ݒ�<��<U��<@��<$��<G��<&��<`   `    ��<U��<t��<I��<@��<S��<R��<:��<t��<2��<���<%��<���<%��<���<2��<t��<:��<R��<S��<@��<I��<t��<U��<`   `   7��<F��<C��<4��<��<��<:��<��<1��<+��< ��</��<��</��< ��<+��<1��<��<:��<��<��<4��<C��<F��<`   `   ؒ�< ��<!��<#��<��<>��<��<В�<'��<H��<A��<��<��<��<A��<H��<'��<В�<��<>��<��<#��<!��< ��<`   `   ��<��<A��<A��<#��<R��<���<��<P��<5��<*��<��<��<��<*��<5��<P��<��<���<R��<#��<A��<A��<��<`   `   0��<=��<:��<^��<A��<��<��<$��<F��<��<8��<��<&��<��<8��<��<F��<$��<��<��<A��<^��<:��<=��<`   `   >��<��<���<��<?��<��<!��<\��<@��<��<!��<��<���<��<!��<��<@��<\��<!��<��<?��<��<���<��<`   `   \��<*��<��<В�<��<I��<-��<I��<(��<+��<��<0��<2��<0��<��<+��<(��<I��<-��<I��<��<В�<��<*��<`   `   H��<��<W��<��<5��<Q��<	��<@��<��<7��<��</��<X��</��<��<7��<��<@��<	��<Q��<5��<��<W��<��<`   `   a��<��<D��<��<��<%��<���<H��<��<+��<���<��<?��<��<���<+��<��<H��<���<%��<��<��<D��<��<`   `   ���< ��<��<��<���<0��<��</��<��<(��<��<��<F��<��<��<(��<��</��<��<0��<���<��<��< ��<`   `   t��< ��<&��<3��<4��<Z��<+��<	��<���<��<&��<*��<��<*��<&��<��<���<	��<+��<Z��<4��<3��<&��< ��<`   `   0��<7��<;��<9��<0��<��<��<��</��<$��<��<��<��<��<��<$��</��<��<��<��<0��<9��<;��<7��<`   `   ���<��<��<&��<��<��<7��<,��<1��<9��<3��<7��<0��<7��<3��<9��<1��<,��<7��<��<��<&��<��<��<`   `   #��<��<��<>��<%��< ��<O��<)��<���<��<>��<W��<W��<W��<>��<��<���<)��<O��< ��<%��<>��<��<��<`   `   ��<8��<4��<5��<=��<'��<!��<��<:��<J��<��<��<��<��<��<J��<:��<��<!��<'��<=��<5��<4��<8��<`   `   ���<#��<��<��<N��<<��<)��<��<.��<a��<��<ؒ�<��<ؒ�<��<a��<.��<��<)��<<��<N��<��<��<#��<`   `   ���<4��<
��<��<'��<��<@��<.��<Ւ�<��<E��<;��<|��<;��<E��<��<Ւ�<.��<@��<��<'��<��<
��<4��<`   `   V��<��<���<`��<R��<��<��<M��<��<��<p��<%��<��<%��<p��<��<��<M��<��<��<R��<`��<���<��<`   `   N��<���<��<h��<~��<V��<���<��<���<;��<j��<��<��<��<j��<;��<���<��<���<V��<~��<h��<��<���<`   `   9��<��<F��<��<��<>��<D��<N��<��<?��<B��<2��<F��<2��<B��<?��<��<N��<D��<>��<��<��<F��<��<`   `   (��<��<C��<��<��<��<8��<`��<3��</��<��<A��<H��<A��<��</��<3��<`��<8��<��<��<��<C��<��<`   `   ��<��<7��<$��<T��<6��<���<��<4��<��<��<X��<K��<X��<��<��<4��<��<���<6��<T��<$��<7��<��<`   `   ��<3��<>��<���<��<��<��<��<1��<��<���<A��<��<A��<���<��<1��<��<��<��<��<���<>��<3��<`   `   ���<<��<.��<��<%��<ݒ�<��<U��<@��<$��<G��<&��<ے�<&��<G��<$��<@��<U��<��<ݒ�<%��<��<.��<<��<`   `   ���<%��<���<2��<t��<:��<R��<S��<@��<I��<t��<U��< ��<U��<t��<I��<@��<S��<R��<:��<t��<2��<���<%��<`   `   ��</��< ��<+��<1��<��<:��<��<��<4��<C��<F��<7��<F��<C��<4��<��<��<:��<��<1��<+��< ��</��<`   `   ��<��<A��<H��<'��<В�<��<>��<��<#��<!��< ��<ؒ�< ��<!��<#��<��<>��<��<В�<'��<H��<A��<��<`   `   ��<��<*��<5��<P��<��<���<R��<#��<A��<A��<��<��<��<A��<A��<#��<R��<���<��<P��<5��<*��<��<`   `   &��<��<8��<��<F��<$��<��<��<A��<^��<:��<=��<0��<=��<:��<^��<A��<��<��<$��<F��<��<8��<��<`   `   ���<��<!��<��<@��<\��<!��<��<?��<��<���<��<>��<��<���<��<?��<��<!��<\��<@��<��<!��<��<`   `   2��<0��<��<+��<(��<I��<-��<I��<��<В�<��<*��<\��<*��<��<В�<��<I��<-��<I��<(��<+��<��<0��<`   `   ���<ٔ�<���<���<���<ޔ�<Ք�<̔�<���<���<��<Ԕ�<���<Ԕ�<��<���<���<̔�<Ք�<ޔ�<���<���<���<ٔ�<`   `   ���<���<���<��<��<	��<��<��<��<
��<*��<Ք�<��<Ք�<*��<
��<��<��<��<	��<��<��<���<���<`   `   Ҕ�<��<���<���< ��<��<Ӕ�< ��<���<���<��<���<��<���<��<���<���< ��<Ӕ�<��< ��<���<���<��<`   `   ϔ�<���<��<���<��<��<��<��<���<Ĕ�<��<���<Ӕ�<���<��<Ĕ�<���<��<��<��<��<���<��<���<`   `   ���<��<ǔ�<��<��<��<ה�<֔�<��<���<��<��< ��<��<��<���<��<֔�<ה�<��<��<��<ǔ�<��<`   `   ۔�<˔�<���<��<۔�<��<��<��<��<Ҕ�<��<ڔ�<��<ڔ�<��<Ҕ�<��<��<��<��<۔�<��<���<˔�<`   `   ���<��<��<֔�<��<���<��<��<Ӕ�<���<��<��<���<��<��<���<Ӕ�<��<��<���<��<֔�<��<��<`   `   Ô�<	��<��<Ȕ�<��<��<���<ɔ�<���<Ȕ�<��<��<���<��<��<Ȕ�<���<ɔ�<���<��<��<Ȕ�<��<	��<`   `   ��<���<���<��<�<��<��<��<��<ɔ�<��<���<���<���<��<ɔ�<��<��<��<��<�<��<���<���<`   `   F��<ޔ�<��<2��<��<���<��<Д�<Δ�<��<���<��<��<��<���<��<Δ�<Д�<��<���<��<2��<��<ޔ�<`   `   ��<���<���<��<3��<��<���<ϔ�<���< ��<��<��<5��<��<��< ��<���<ϔ�<���<��<3��<��<���<���<`   `   ��<��<���<Ҕ�<��<��<��<���<Ȕ�<͔�<��<Ӕ�<��<Ӕ�<��<͔�<Ȕ�<���<��<��<��<Ҕ�<���<��<`   `   ��<;��<��<��<��<ޔ�<���<ܔ�<ʔ�<���<��<��<���<��<��<���<ʔ�<ܔ�<���<ޔ�<��<��<��<;��<`   `   ���<Ք�<���<��<��<���<��<ϔ�<��<ٔ�<���<��<���<��<���<ٔ�<��<ϔ�<��<���<��<��<���<Ք�<`   `   ���<��<��<5��<��<��<��<��<2��<��<���<��<��<��<���<��<2��<��<��<��<��<5��<��<��<`   `   ǔ�<S��<I��<��<���<��<4��<���<��<��<���<���<��<���<���<��<��<���<4��<��<���<��<I��<S��<`   `   є�<��<��<���<ޔ�<Δ�< ��<��<��<���<��<��<���<��<��<���<��<��< ��<Δ�<ޔ�<���<��<��<`   `   %��<���<���<���< ��<���<є�<��<͔�<��<��<��<ߔ�<��<��<��<͔�<��<є�<���< ��<���<���<���<`   `   ���<֔�<۔�<��<��<���<Ô�<��<���<֔�<��<��<��<��<��<֔�<���<��<Ô�<���<��<��<۔�<֔�<`   `   E��<ϔ�<���<��<є�<+��<��<��<��<̔�<ה�<��<��<��<ה�<̔�<��<��<��<+��<є�<��<���<ϔ�<`   `   &��<���<��<���<���<C��<��<��<��<���<̔�<��<	��<��<̔�<���<��<��<��<C��<���<���<��<���<`   `   ��<��<Ô�<���<���<ה�<��<���<Δ�<Ŕ�< ��<���<��<���< ��<Ŕ�<Δ�<���<��<ה�<���<���<Ô�<��<`   `   ���<��<��</��<��<���<��<Ԕ�<ؔ�<��<��<ٔ�<���<ٔ�<��<��<ؔ�<Ԕ�<��<���<��</��<��<��<`   `   ܔ�<��<��<!��< ��<���<��<���<���<���<Ӕ�<Ԕ�<���<Ԕ�<Ӕ�<���<���<���<��<���< ��<!��<��<��<`   `   ���<Ԕ�<��<���<���<̔�<Ք�<ޔ�<���<���<���<ٔ�<���<ٔ�<���<���<���<ޔ�<Ք�<̔�<���<���<��<Ԕ�<`   `   ��<Ք�<*��<
��<��<��<��<	��<��<��<���<���<���<���<���<��<��<	��<��<��<��<
��<*��<Ք�<`   `   ��<���<��<���<���< ��<Ӕ�<��< ��<���<���<��<Ҕ�<��<���<���< ��<��<Ӕ�< ��<���<���<��<���<`   `   Ӕ�<���<��<Ĕ�<���<��<��<��<��<���<��<���<ϔ�<���<��<���<��<��<��<��<���<Ĕ�<��<���<`   `    ��<��<��<���<��<֔�<ה�<��<��<��<ǔ�<��<���<��<ǔ�<��<��<��<ה�<֔�<��<���<��<��<`   `   ��<ڔ�<��<Ҕ�<��<��<��<��<۔�<��<���<˔�<۔�<˔�<���<��<۔�<��<��<��<��<Ҕ�<��<ڔ�<`   `   ���<��<��<���<Ӕ�<��<��<���<��<֔�<��<��<���<��<��<֔�<��<���<��<��<Ӕ�<���<��<��<`   `   ���<��<��<Ȕ�<���<ɔ�<���<��<��<Ȕ�<��<	��<Ô�<	��<��<Ȕ�<��<��<���<ɔ�<���<Ȕ�<��<��<`   `   ���<���<��<ɔ�<��<��<��<��<�<��<���<���<��<���<���<��<�<��<��<��<��<ɔ�<��<���<`   `   ��<��<���<��<Δ�<Д�<��<���<��<2��<��<ޔ�<F��<ޔ�<��<2��<��<���<��<Д�<Δ�<��<���<��<`   `   5��<��<��< ��<���<ϔ�<���<��<3��<��<���<���<��<���<���<��<3��<��<���<ϔ�<���< ��<��<��<`   `   ��<Ӕ�<��<͔�<Ȕ�<���<��<��<��<Ҕ�<���<��<��<��<���<Ҕ�<��<��<��<���<Ȕ�<͔�<��<Ӕ�<`   `   ���<��<��<���<ʔ�<ܔ�<���<ޔ�<��<��<��<;��<��<;��<��<��<��<ޔ�<���<ܔ�<ʔ�<���<��<��<`   `   ���<��<���<ٔ�<��<ϔ�<��<���<��<��<���<Ք�<���<Ք�<���<��<��<���<��<ϔ�<��<ٔ�<���<��<`   `   ��<��<���<��<2��<��<��<��<��<5��<��<��<���<��<��<5��<��<��<��<��<2��<��<���<��<`   `   ��<���<���<��<��<���<4��<��<���<��<I��<S��<ǔ�<S��<I��<��<���<��<4��<���<��<��<���<���<`   `   ���<��<��<���<��<��< ��<Δ�<ޔ�<���<��<��<є�<��<��<���<ޔ�<Δ�< ��<��<��<���<��<��<`   `   ߔ�<��<��<��<͔�<��<є�<���< ��<���<���<���<%��<���<���<���< ��<���<є�<��<͔�<��<��<��<`   `   ��<��<��<֔�<���<��<Ô�<���<��<��<۔�<֔�<���<֔�<۔�<��<��<���<Ô�<��<���<֔�<��<��<`   `   ��<��<ה�<̔�<��<��<��<+��<є�<��<���<ϔ�<E��<ϔ�<���<��<є�<+��<��<��<��<̔�<ה�<��<`   `   	��<��<̔�<���<��<��<��<C��<���<���<��<���<&��<���<��<���<���<C��<��<��<��<���<̔�<��<`   `   ��<���< ��<Ŕ�<Δ�<���<��<ה�<���<���<Ô�<��<��<��<Ô�<���<���<ה�<��<���<Δ�<Ŕ�< ��<���<`   `   ���<ٔ�<��<��<ؔ�<Ԕ�<��<���<��</��<��<��<���<��<��</��<��<���<��<Ԕ�<ؔ�<��<��<ٔ�<`   `   ���<Ԕ�<Ӕ�<���<���<���<��<���< ��<!��<��<��<ܔ�<��<��<!��< ��<���<��<���<���<���<Ӕ�<Ԕ�<`   `   ���<Ȗ�<���<���<��<ϖ�<��<���<ɖ�<���<���<ʖ�<Ӗ�<ʖ�<���<���<ɖ�<���<��<ϖ�<��<���<���<Ȗ�<`   `   ���<��<���<���<Ŗ�<���<ݖ�<���<ϖ�<���<���<��<���<��<���<���<ϖ�<���<ݖ�<���<Ŗ�<���<���<��<`   `   ���<���<|��<���<���<���<���<z��<���<���<Ŗ�<��<���<��<Ŗ�<���<���<z��<���<���<���<���<|��<���<`   `   ~��<���<���<���<���<Ö�<ۖ�<���<Ζ�<���<���<Ֆ�<���<Ֆ�<���<���<Ζ�<���<ۖ�<Ö�<���<���<���<���<`   `   Ӗ�<Ж�<��<Ö�<���<ܖ�<˖�<���<ϖ�<���<���<���<Ö�<���<���<���<ϖ�<���<˖�<ܖ�<���<Ö�<��<Ж�<`   `   ֖�<Ɩ�<Ԗ�<ۖ�<���<���<���<���<ϖ�<���<Ȗ�<�<��<�<Ȗ�<���<ϖ�<���<���<���<���<ۖ�<Ԗ�<Ɩ�<`   `   ���<���<���<��<Җ�<|��<���<ܖ�<˖�<��<ۖ�<���<���<���<ۖ�<��<˖�<ܖ�<���<|��<Җ�<��<���<���<`   `   Ֆ�<��<���<���<̖�<���<ϖ�<̖�<���<ݖ�<���<f��<Җ�<f��<���<ݖ�<���<̖�<ϖ�<���<̖�<���<���<��<`   `   ���<Ɩ�<���<���<���<ߖ�<���<���<���<ǖ�<���<���<'��<���<���<ǖ�<���<���<���<ߖ�<���<���<���<Ɩ�<`   `   T��<���<֖�<���<͖�<���<���<��<ז�<і�<і�<���<Ŗ�<���<і�<і�<ז�<��<���<���<͖�<���<֖�<���<`   `   Ɩ�<��<��<���<Ė�<z��<Ȗ�<��<���<���<і�<���<^��<���<і�<���<���<��<Ȗ�<z��<Ė�<���<��<��<`   `   ���<��<ז�<���<Ȗ�<���<Ӗ�<���<���<���<���<Ӗ�<���<Ӗ�<���<���<���<���<Ӗ�<���<Ȗ�<���<ז�<��<`   `   X��<���<Ԗ�<ۖ�<ז�<��<Ȗ�<���<��<��<���<ǖ�<ږ�<ǖ�<���<��<��<���<Ȗ�<��<ז�<ۖ�<Ԗ�<���<`   `   ���<���<ݖ�<���<���<̖�<ܖ�<�<ޖ�<ɖ�<���<���<Ȗ�<���<���<ɖ�<ޖ�<�<ܖ�<̖�<���<���<ݖ�<���<`   `    ��<Җ�<���<���<���<͖�<ϖ�<���<c��<���<і�<���<̖�<���<і�<���<c��<���<ϖ�<͖�<���<���<���<Җ�<`   `   ݖ�<}��<���<ޖ�<ϖ�<���<���<���<���<��<���<���<���<���<���<��<���<���<���<���<ϖ�<ޖ�<���<}��<`   `   S��<˖�<֖�<��<̖�<���<���<͖�<̖�<̖�<v��<���<ܖ�<���<v��<̖�<̖�<͖�<���<���<̖�<��<֖�<˖�<`   `   Ԗ�<�<��<���<��<	��<і�<���<���<Ӗ�<���<���<ߖ�<���<���<Ӗ�<���<���<і�<	��<��<���<��<�<`   `   l��<���<��<m��<֖�<��<���<Ɩ�<���<���<ϖ�<���<���<���<ϖ�<���<���<Ɩ�<���<��<֖�<m��<��<���<`   `   ���<ږ�<��<���<Җ�<���<m��<Ֆ�<���<Ζ�<֖�<���<���<���<֖�<Ζ�<���<Ֆ�<m��<���<Җ�<���<��<ږ�<`   `   ���<Ɩ�<���<��<��<v��<���<ǖ�<���<�<ޖ�<���<���<���<ޖ�<�<���<ǖ�<���<v��<��<��<���<Ɩ�<`   `   o��<Ֆ�<���<˖�<��<���<��<Ֆ�<Ŗ�<і�<ɖ�<���<���<���<ɖ�<і�<Ŗ�<Ֆ�<��<���<��<˖�<���<Ֆ�<`   `   ���<��<���<���<���<���<Ԗ�<Ŗ�<ؖ�<���<���<���<���<���<���<���<ؖ�<Ŗ�<Ԗ�<���<���<���<���<��<`   `   ٖ�<ݖ�<���<���<���<���<���<���<��<���<���<ɖ�<���<ɖ�<���<���<��<���<���<���<���<���<���<ݖ�<`   `   Ӗ�<ʖ�<���<���<ɖ�<���<��<ϖ�<��<���<���<Ȗ�<���<Ȗ�<���<���<��<ϖ�<��<���<ɖ�<���<���<ʖ�<`   `   ���<��<���<���<ϖ�<���<ݖ�<���<Ŗ�<���<���<��<���<��<���<���<Ŗ�<���<ݖ�<���<ϖ�<���<���<��<`   `   ���<��<Ŗ�<���<���<z��<���<���<���<���<|��<���<���<���<|��<���<���<���<���<z��<���<���<Ŗ�<��<`   `   ���<Ֆ�<���<���<Ζ�<���<ۖ�<Ö�<���<���<���<���<~��<���<���<���<���<Ö�<ۖ�<���<Ζ�<���<���<Ֆ�<`   `   Ö�<���<���<���<ϖ�<���<˖�<ܖ�<���<Ö�<��<Ж�<Ӗ�<Ж�<��<Ö�<���<ܖ�<˖�<���<ϖ�<���<���<���<`   `   ��<�<Ȗ�<���<ϖ�<���<���<���<���<ۖ�<Ԗ�<Ɩ�<֖�<Ɩ�<Ԗ�<ۖ�<���<���<���<���<ϖ�<���<Ȗ�<�<`   `   ���<���<ۖ�<��<˖�<ܖ�<���<|��<Җ�<��<���<���<���<���<���<��<Җ�<|��<���<ܖ�<˖�<��<ۖ�<���<`   `   Җ�<f��<���<ݖ�<���<̖�<ϖ�<���<̖�<���<���<��<Ֆ�<��<���<���<̖�<���<ϖ�<̖�<���<ݖ�<���<f��<`   `   '��<���<���<ǖ�<���<���<���<ߖ�<���<���<���<Ɩ�<���<Ɩ�<���<���<���<ߖ�<���<���<���<ǖ�<���<���<`   `   Ŗ�<���<і�<і�<ז�<��<���<���<͖�<���<֖�<���<T��<���<֖�<���<͖�<���<���<��<ז�<і�<і�<���<`   `   ^��<���<і�<���<���<��<Ȗ�<z��<Ė�<���<��<��<Ɩ�<��<��<���<Ė�<z��<Ȗ�<��<���<���<і�<���<`   `   ���<Ӗ�<���<���<���<���<Ӗ�<���<Ȗ�<���<ז�<��<���<��<ז�<���<Ȗ�<���<Ӗ�<���<���<���<���<Ӗ�<`   `   ږ�<ǖ�<���<��<��<���<Ȗ�<��<ז�<ۖ�<Ԗ�<���<X��<���<Ԗ�<ۖ�<ז�<��<Ȗ�<���<��<��<���<ǖ�<`   `   Ȗ�<���<���<ɖ�<ޖ�<�<ܖ�<̖�<���<���<ݖ�<���<���<���<ݖ�<���<���<̖�<ܖ�<�<ޖ�<ɖ�<���<���<`   `   ̖�<���<і�<���<c��<���<ϖ�<͖�<���<���<���<Җ�< ��<Җ�<���<���<���<͖�<ϖ�<���<c��<���<і�<���<`   `   ���<���<���<��<���<���<���<���<ϖ�<ޖ�<���<}��<ݖ�<}��<���<ޖ�<ϖ�<���<���<���<���<��<���<���<`   `   ܖ�<���<v��<̖�<̖�<͖�<���<���<̖�<��<֖�<˖�<S��<˖�<֖�<��<̖�<���<���<͖�<̖�<̖�<v��<���<`   `   ߖ�<���<���<Ӗ�<���<���<і�<	��<��<���<��<�<Ԗ�<�<��<���<��<	��<і�<���<���<Ӗ�<���<���<`   `   ���<���<ϖ�<���<���<Ɩ�<���<��<֖�<m��<��<���<l��<���<��<m��<֖�<��<���<Ɩ�<���<���<ϖ�<���<`   `   ���<���<֖�<Ζ�<���<Ֆ�<m��<���<Җ�<���<��<ږ�<���<ږ�<��<���<Җ�<���<m��<Ֆ�<���<Ζ�<֖�<���<`   `   ���<���<ޖ�<�<���<ǖ�<���<v��<��<��<���<Ɩ�<���<Ɩ�<���<��<��<v��<���<ǖ�<���<�<ޖ�<���<`   `   ���<���<ɖ�<і�<Ŗ�<Ֆ�<��<���<��<˖�<���<Ֆ�<o��<Ֆ�<���<˖�<��<���<��<Ֆ�<Ŗ�<і�<ɖ�<���<`   `   ���<���<���<���<ؖ�<Ŗ�<Ԗ�<���<���<���<���<��<���<��<���<���<���<���<Ԗ�<Ŗ�<ؖ�<���<���<���<`   `   ���<ɖ�<���<���<��<���<���<���<���<���<���<ݖ�<ٖ�<ݖ�<���<���<���<���<���<���<��<���<���<ɖ�<`   `   ���<u��<���<���<���<e��<���<���<���<��<ט�<���<���<���<ט�<��<���<���<���<e��<���<���<���<u��<`   `   ���<p��<���<���<���<h��<���<z��<���<���<���<���<L��<���<���<���<���<z��<���<h��<���<���<���<p��<`   `   ���<���<���<���<���<���<ژ�<���<���<���<b��<���<k��<���<b��<���<���<���<ژ�<���<���<���<���<���<`   `   Ԙ�<���<���<���<���<s��<���<���<���<ј�<���<���<���<���<���<ј�<���<���<���<s��<���<���<���<���<`   `   }��<_��<���<���<���<���<l��<���<���<���<���<���<��<���<���<���<���<���<l��<���<���<���<���<_��<`   `   }��<���<���<^��<���<��<���<���<|��<{��<���<���<���<���<���<{��<|��<���<���<��<���<^��<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<r��<���<ݘ�<���<l��<ɘ�<���<���<���<���<���<���<���<���<���<���<���<ɘ�<l��<���<ݘ�<���<r��<`   `   Ø�<���<���<ј�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<ј�<���<���<`   `   ǘ�<���<���<���<���<ט�<r��<s��<���<���<���<���<���<���<���<���<���<s��<r��<ט�<���<���<���<���<`   `   ���<���<���<���<���<��<���<���<���<���<���<���<���<���<���<���<���<���<���<��<���<���<���<���<`   `   Ř�<~��<���<���<y��<���<���<[��<���<���<���<���<���<���<���<���<���<[��<���<���<y��<���<���<~��<`   `   �<e��<���<���<���<���<���<���<���<���<v��<���<���<���<v��<���<���<���<���<���<���<���<���<e��<`   `   ��<���<˘�<���<���<Ę�<���<��<g��<z��<���<���<���<���<���<z��<g��<��<���<Ę�<���<���<˘�<���<`   `   ǘ�<���<ݘ�<���<Ș�<���<g��<��<���<���<ݘ�<���<���<���<ݘ�<���<���<��<g��<���<Ș�<���<ݘ�<���<`   `   ���<v��<���<���<���<���<p��<͘�<՘�<���<���<���<���<���<���<���<՘�<͘�<p��<���<���<���<���<v��<`   `   ͘�<���<���<���<���<���<���<���<���<v��<���<�<t��<�<���<v��<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<l��<���<���<���<���<���<���<���<]��<���<���<���<���<���<���<���<l��<���<���<���<`   `   ���<ʘ�<И�<���<���<���<���<���<ޘ�<���<q��<���<x��<���<q��<���<ޘ�<���<���<���<���<���<И�<ʘ�<`   `   Ҙ�<Θ�<���<���<���<���<ј�<���<{��<k��<c��<���<���<���<c��<k��<{��<���<ј�<���<���<���<���<Θ�<`   `   ���<���<���<���<���<���<ޘ�<���<}��<���<���<���<���<���<���<���<}��<���<ޘ�<���<���<���<���<���<`   `   �<՘�<Ә�<���<Ř�<���<���<���<���<���<n��<���<̘�<���<n��<���<���<���<���<���<Ř�<���<Ә�<՘�<`   `   ؘ�<���<���<t��<���<���<^��<���<���<k��<���<���<���<���<���<k��<���<���<^��<���<���<t��<���<���<`   `   ���<���<���<���<���<֘�<���<���<���<���<Ԙ�<���<i��<���<Ԙ�<���<���<���<���<֘�<���<���<���<���<`   `   ���<���<ט�<��<���<���<���<e��<���<���<���<u��<���<u��<���<���<���<e��<���<���<���<��<ט�<���<`   `   L��<���<���<���<���<z��<���<h��<���<���<���<p��<���<p��<���<���<���<h��<���<z��<���<���<���<���<`   `   k��<���<b��<���<���<���<ژ�<���<���<���<���<���<���<���<���<���<���<���<ژ�<���<���<���<b��<���<`   `   ���<���<���<ј�<���<���<���<s��<���<���<���<���<Ԙ�<���<���<���<���<s��<���<���<���<ј�<���<���<`   `   ��<���<���<���<���<���<l��<���<���<���<���<_��<}��<_��<���<���<���<���<l��<���<���<���<���<���<`   `   ���<���<���<{��<|��<���<���<��<���<^��<���<���<}��<���<���<^��<���<��<���<���<|��<{��<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<���<���<ɘ�<l��<���<ݘ�<���<r��<���<r��<���<ݘ�<���<l��<ɘ�<���<���<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<ј�<���<���<Ø�<���<���<ј�<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<���<s��<r��<ט�<���<���<���<���<ǘ�<���<���<���<���<ט�<r��<s��<���<���<���<���<`   `   ���<���<���<���<���<���<���<��<���<���<���<���<���<���<���<���<���<��<���<���<���<���<���<���<`   `   ���<���<���<���<���<[��<���<���<y��<���<���<~��<Ř�<~��<���<���<y��<���<���<[��<���<���<���<���<`   `   ���<���<v��<���<���<���<���<���<���<���<���<e��<�<e��<���<���<���<���<���<���<���<���<v��<���<`   `   ���<���<���<z��<g��<��<���<Ę�<���<���<˘�<���<��<���<˘�<���<���<Ę�<���<��<g��<z��<���<���<`   `   ���<���<ݘ�<���<���<��<g��<���<Ș�<���<ݘ�<���<ǘ�<���<ݘ�<���<Ș�<���<g��<��<���<���<ݘ�<���<`   `   ���<���<���<���<՘�<͘�<p��<���<���<���<���<v��<���<v��<���<���<���<���<p��<͘�<՘�<���<���<���<`   `   t��<�<���<v��<���<���<���<���<���<���<���<���<͘�<���<���<���<���<���<���<���<���<v��<���<�<`   `   ]��<���<���<���<���<���<���<���<l��<���<���<���<���<���<���<���<l��<���<���<���<���<���<���<���<`   `   x��<���<q��<���<ޘ�<���<���<���<���<���<И�<ʘ�<���<ʘ�<И�<���<���<���<���<���<ޘ�<���<q��<���<`   `   ���<���<c��<k��<{��<���<ј�<���<���<���<���<Θ�<Ҙ�<Θ�<���<���<���<���<ј�<���<{��<k��<c��<���<`   `   ���<���<���<���<}��<���<ޘ�<���<���<���<���<���<���<���<���<���<���<���<ޘ�<���<}��<���<���<���<`   `   ̘�<���<n��<���<���<���<���<���<Ř�<���<Ә�<՘�<�<՘�<Ә�<���<Ř�<���<���<���<���<���<n��<���<`   `   ���<���<���<k��<���<���<^��<���<���<t��<���<���<ؘ�<���<���<t��<���<���<^��<���<���<k��<���<���<`   `   i��<���<Ԙ�<���<���<���<���<֘�<���<���<���<���<���<���<���<���<���<֘�<���<���<���<���<Ԙ�<���<`   `   ��<k��<b��<i��<|��<���<X��<p��<T��<g��<���<���<���<���<���<g��<T��<p��<X��<���<|��<i��<b��<k��<`   `   ���<V��<���<_��<���<���<a��<���<��<���<���<���<���<���<���<���<��<���<a��<���<���<_��<���<V��<`   `   J��<E��<���<.��<q��<���<s��<���<���<���<���<���<���<���<���<���<���<���<s��<���<q��<.��<���<E��<`   `   ���<w��<y��<N��<���<���<P��<s��<,��<w��<���<���<���<���<���<w��<,��<s��<P��<���<���<N��<y��<w��<`   `   ���<j��<���<���<���<a��<���<���<[��<���<���<���<���<���<���<���<[��<���<���<a��<���<���<���<j��<`   `   ~��<���<���<���<���<_��<���<���<���<���<���<���<g��<���<���<���<���<���<���<_��<���<���<���<���<`   `   ���<���<���<i��<���<���<[��<S��<ƚ�<u��<J��<���<f��<���<J��<u��<ƚ�<S��<[��<���<���<i��<���<���<`   `   l��<u��<���<r��<{��<���<^��<c��<���<c��<p��<���<U��<���<p��<c��<���<c��<^��<���<{��<r��<���<u��<`   `   ���<���<���<���<k��<}��<���<���<���<���<���<���<@��<���<���<���<���<���<���<}��<k��<���<���<���<`   `   ˚�<���<���<���<r��<���<���<���<���<���<y��<���<���<���<y��<���<���<���<���<���<r��<���<���<���<`   `   ~��<P��<���<Ś�<���<���<���<���<���<���<|��<���<���<���<|��<���<���<���<���<���<���<Ś�<���<P��<`   `   ��<���<���<ƚ�<���<���<���<Ț�<���<���<���<q��<3��<q��<���<���<���<Ț�<���<���<���<ƚ�<���<���<`   `   ��<ؚ�<���<l��<���<u��<���<Ś�<k��<���<���<���<a��<���<���<���<k��<Ś�<���<u��<���<l��<���<ؚ�<`   `   \��<[��<���<���<���<���<~��<���<|��<���<���<���<���<���<���<���<|��<���<~��<���<���<���<���<[��<`   `   {��<���<���<���<���<���<���<���<���<���<:��<c��<���<c��<:��<���<���<���<���<���<���<���<���<���<`   `   ˚�<��<՚�<z��<o��<���<���<u��<��<q��<K��<}��<���<}��<K��<q��<��<u��<���<���<o��<z��<՚�<��<`   `   e��<Κ�<���<���<���<͚�<ښ�<u��<e��<���<���<z��<t��<z��<���<���<e��<u��<ښ�<͚�<���<���<���<Κ�<`   `   ���<���<8��<���<���<q��<���<���<���<y��<���<j��<f��<j��<���<y��<���<���<���<q��<���<���<8��<���<`   `   ���<���<S��<��<�<V��<{��<r��<���<a��<~��<���<���<���<~��<a��<���<r��<{��<V��<�<��<S��<���<`   `   ���<���<���<��<���<���<���<g��<���<���<���<���<V��<���<���<���<���<g��<���<���<���<��<���<���<`   `   ���<���<���<���<S��<���<���<���<���<���<��<w��< ��<w��<��<���<���<���<���<���<S��<���<���<���<`   `   ���<e��<���<���<z��<z��<p��<���<���<x��<\��<���<q��<���<\��<x��<���<���<p��<z��<z��<���<���<e��<`   `   ���<^��<���<Ԛ�<���<���<���<���<r��<���<���<j��<h��<j��<���<���<r��<���<���<���<���<Ԛ�<���<^��<`   `   ���<x��<���<���<y��<���<���<К�<x��<���<x��<E��<���<E��<x��<���<x��<К�<���<���<y��<���<���<x��<`   `   ���<���<���<g��<T��<p��<X��<���<|��<i��<b��<k��<��<k��<b��<i��<|��<���<X��<p��<T��<g��<���<���<`   `   ���<���<���<���<��<���<a��<���<���<_��<���<V��<���<V��<���<_��<���<���<a��<���<��<���<���<���<`   `   ���<���<���<���<���<���<s��<���<q��<.��<���<E��<J��<E��<���<.��<q��<���<s��<���<���<���<���<���<`   `   ���<���<���<w��<,��<s��<P��<���<���<N��<y��<w��<���<w��<y��<N��<���<���<P��<s��<,��<w��<���<���<`   `   ���<���<���<���<[��<���<���<a��<���<���<���<j��<���<j��<���<���<���<a��<���<���<[��<���<���<���<`   `   g��<���<���<���<���<���<���<_��<���<���<���<���<~��<���<���<���<���<_��<���<���<���<���<���<���<`   `   f��<���<J��<u��<ƚ�<S��<[��<���<���<i��<���<���<���<���<���<i��<���<���<[��<S��<ƚ�<u��<J��<���<`   `   U��<���<p��<c��<���<c��<^��<���<{��<r��<���<u��<l��<u��<���<r��<{��<���<^��<c��<���<c��<p��<���<`   `   @��<���<���<���<���<���<���<}��<k��<���<���<���<���<���<���<���<k��<}��<���<���<���<���<���<���<`   `   ���<���<y��<���<���<���<���<���<r��<���<���<���<ʚ�<���<���<���<r��<���<���<���<���<���<y��<���<`   `   ���<���<|��<���<���<���<���<���<���<Ś�<���<P��<~��<P��<���<Ś�<���<���<���<���<���<���<|��<���<`   `   3��<q��<���<���<���<Ț�<���<���<���<ƚ�<���<���<��<���<���<ƚ�<���<���<���<Ț�<���<���<���<q��<`   `   a��<���<���<���<k��<Ś�<���<u��<���<l��<���<ؚ�<��<ؚ�<���<l��<���<u��<���<Ś�<k��<���<���<���<`   `   ���<���<���<���<|��<���<~��<���<���<���<���<[��<\��<[��<���<���<���<���<~��<���<|��<���<���<���<`   `   ���<c��<:��<���<���<���<���<���<���<���<���<���<{��<���<���<���<���<���<���<���<���<���<:��<c��<`   `   ���<}��<K��<q��<��<u��<���<���<o��<z��<՚�<��<˚�<��<՚�<z��<o��<���<���<u��<��<q��<K��<}��<`   `   t��<z��<���<���<e��<u��<ښ�<͚�<���<���<���<Κ�<e��<Κ�<���<���<���<͚�<ښ�<u��<e��<���<���<z��<`   `   f��<j��<���<y��<���<���<���<q��<���<���<8��<���<���<���<8��<���<���<q��<���<���<���<y��<���<j��<`   `   ���<���<~��<a��<���<r��<{��<V��<�<��<S��<���<���<���<S��<��<�<V��<{��<r��<���<a��<~��<���<`   `   V��<���<���<���<���<g��<���<���<���<��<���<���<���<���<���<��<���<���<���<g��<���<���<���<���<`   `    ��<w��<��<���<���<���<���<���<S��<���<���<���<���<���<���<���<S��<���<���<���<���<���<��<w��<`   `   q��<���<\��<x��<���<���<p��<z��<z��<���<���<e��<���<e��<���<���<z��<z��<p��<���<���<x��<\��<���<`   `   h��<j��<���<���<r��<���<���<���<���<Ԛ�<���<^��<���<^��<���<Ԛ�<���<���<���<���<r��<���<���<j��<`   `   ���<E��<x��<���<x��<К�<���<���<y��<���<���<x��<���<x��<���<���<y��<���<���<К�<x��<���<x��<E��<`   `   :��<v��<w��<q��<t��<k��<���<���<���<���<R��<d��<r��<d��<R��<���<���<���<���<k��<t��<q��<w��<v��<`   `   o��<���<���<���<���<l��<���<���<���<���<���<o��<���<o��<���<���<���<���<���<l��<���<���<���<���<`   `   ���<v��<z��<���<^��<?��<E��<���<���<���<���<���<���<���<���<���<���<���<E��<?��<^��<���<z��<v��<`   `   R��<e��<���<���<b��<���<���<���<���<x��<|��<t��<f��<t��<|��<x��<���<���<���<���<b��<���<���<e��<`   `   z��<���<s��<k��<X��<���<���<r��<���<~��<`��<���<���<���<`��<~��<���<r��<���<���<X��<k��<s��<���<`   `   l��<S��<F��<���<`��<2��<���<N��<0��<��<���<���<���<���<���<��<0��<N��<���<2��<`��<���<F��<S��<`   `   i��<O��<`��<���<���<��<���<���<Q��<���<���<}��<t��<}��<���<���<Q��<���<���<��<���<���<`��<O��<`   `   ���<���<���<g��<���<���<���<���<q��<���<���<���<���<���<���<���<q��<���<���<���<���<g��<���<���<`   `   D��<x��<���<���<���<���<t��<b��<N��<���<o��<���<���<���<o��<���<N��<b��<t��<���<���<���<���<x��<`   `   T��<���<���<���<���<���<���<���<b��<���<���<l��<���<l��<���<���<b��<���<���<���<���<���<���<���<`   `   ���<��<���<c��<v��<Y��<i��<v��<g��<���<���<s��<���<s��<���<���<g��<v��<i��<Y��<v��<c��<���<��<`   `   ��<���<���<W��<���<���<j��<���<w��<r��<���<���<���<���<���<r��<w��<���<j��<���<���<W��<���<���<`   `   +��<���<���<y��<���<���<���<���<���<}��<a��<���<���<���<a��<}��<���<���<���<���<���<y��<���<���<`   `   Ŝ�<ʜ�<Ȝ�<���<���<���<���<F��<���<���<T��<���<Q��<���<T��<���<���<F��<���<���<���<���<Ȝ�<ʜ�<`   `   ��<���<b��<ڜ�<���<���<��<Y��<���<���<���<���<7��<���<���<���<���<Y��<��<���<���<ڜ�<b��<���<`   `   ���<���<G��<Ĝ�<���<R��<���<u��<���<���<���<���<���<���<���<���<���<u��<���<R��<���<Ĝ�<G��<���<`   `   #��<���<���<Ҝ�<���<Y��<O��<���<���<���<���<L��<���<L��<���<���<���<���<O��<Y��<���<Ҝ�<���<���<`   `   ���<��<���<���<���<ǜ�<���<���<���<���<p��<2��<ݜ�<2��<p��<���<���<���<���<ǜ�<���<���<���<��<`   `   x��<���<���<L��<A��<���<���<���<i��<���<���<9��<���<9��<���<���<i��<���<���<���<A��<L��<���<���<`   `   R��<���<���<f��<x��<���<S��<���<���<���<���<J��<q��<J��<���<���<���<���<S��<���<x��<f��<���<���<`   `   Ԝ�<̜�<М�<���<��<���<*��<���<]��<C��<n��<���<���<���<n��<C��<]��<���<*��<���<��<���<М�<̜�<`   `   Ĝ�<���<j��<i��<͜�<���<���<���<N��<g��<v��<���<S��<���<v��<g��<N��<���<���<���<͜�<i��<j��<���<`   `   ���<���<���<_��<���<{��<���<^��<h��<���<d��<���<l��<���<d��<���<h��<^��<���<{��<���<_��<���<���<`   `   ���<ǜ�<���<���<���<t��<u��<=��<\��<���<G��<���<{��<���<G��<���<\��<=��<u��<t��<���<���<���<ǜ�<`   `   r��<d��<R��<���<���<���<���<k��<t��<q��<w��<v��<:��<v��<w��<q��<t��<k��<���<���<���<���<R��<d��<`   `   ���<o��<���<���<���<���<���<l��<���<���<���<���<o��<���<���<���<���<l��<���<���<���<���<���<o��<`   `   ���<���<���<���<���<���<E��<?��<^��<���<z��<v��<���<v��<z��<���<^��<?��<E��<���<���<���<���<���<`   `   f��<t��<|��<x��<���<���<���<���<b��<���<���<e��<R��<e��<���<���<b��<���<���<���<���<x��<|��<t��<`   `   ���<���<`��<~��<���<r��<���<���<X��<k��<s��<���<z��<���<s��<k��<X��<���<���<r��<���<~��<`��<���<`   `   ���<���<���<��<0��<N��<���<2��<`��<���<F��<S��<l��<S��<F��<���<`��<2��<���<N��<0��<��<���<���<`   `   t��<}��<���<���<Q��<���<���<��<���<���<`��<O��<i��<O��<`��<���<���<��<���<���<Q��<���<���<}��<`   `   ���<���<���<���<q��<���<���<���<���<g��<���<���<���<���<���<g��<���<���<���<���<q��<���<���<���<`   `   ���<���<o��<���<N��<b��<t��<���<���<���<���<x��<D��<x��<���<���<���<���<t��<b��<N��<���<o��<���<`   `   ���<l��<���<���<b��<���<���<���<���<���<���<���<T��<���<���<���<���<���<���<���<b��<���<���<l��<`   `   ���<s��<���<���<g��<v��<i��<Y��<v��<c��<���<��<���<��<���<c��<v��<Y��<i��<v��<g��<���<���<s��<`   `   ���<���<���<r��<w��<���<j��<���<���<W��<���<���<��<���<���<W��<���<���<j��<���<w��<r��<���<���<`   `   ���<���<a��<}��<���<���<���<���<���<y��<���<���<+��<���<���<y��<���<���<���<���<���<}��<a��<���<`   `   Q��<���<T��<���<���<F��<���<���<���<���<Ȝ�<ʜ�<Ŝ�<ʜ�<Ȝ�<���<���<���<���<F��<���<���<T��<���<`   `   7��<���<���<���<���<Y��<��<���<���<ڜ�<b��<���<��<���<b��<ڜ�<���<���<��<Y��<���<���<���<���<`   `   ���<���<���<���<���<u��<���<R��<���<Ĝ�<G��<���<���<���<G��<Ĝ�<���<R��<���<u��<���<���<���<���<`   `   ���<L��<���<���<���<���<O��<Y��<���<Ҝ�<���<���<#��<���<���<Ҝ�<���<Y��<O��<���<���<���<���<L��<`   `   ݜ�<2��<p��<���<���<���<���<ǜ�<���<���<���<��<���<��<���<���<���<ǜ�<���<���<���<���<p��<2��<`   `   ���<9��<���<���<i��<���<���<���<A��<L��<���<���<x��<���<���<L��<A��<���<���<���<i��<���<���<9��<`   `   q��<J��<���<���<���<���<S��<���<x��<f��<���<���<R��<���<���<f��<x��<���<S��<���<���<���<���<J��<`   `   ���<���<n��<C��<]��<���<*��<���<��<���<М�<̜�<Ԝ�<̜�<М�<���<��<���<*��<���<]��<C��<n��<���<`   `   S��<���<v��<g��<N��<���<���<���<͜�<i��<j��<���<Ĝ�<���<j��<i��<͜�<���<���<���<N��<g��<v��<���<`   `   l��<���<d��<���<h��<^��<���<{��<���<_��<���<���<���<���<���<_��<���<{��<���<^��<h��<���<d��<���<`   `   {��<���<G��<���<\��<=��<u��<t��<���<���<���<ǜ�<���<ǜ�<���<���<���<t��<u��<=��<\��<���<G��<���<`   `   ֝�<l��<���<k��<z��<���<���<N��<���<���<���<�<���<�<���<���<���<N��<���<���<z��<k��<���<l��<`   `   I��<j��<*��<Y��<r��<z��<���<D��<=��<���<���<���<���<���<���<���<=��<D��<���<z��<r��<Y��<*��<j��<`   `   ���<���<��<���<���<v��<���<j��<V��<T��<���<~��<���<~��<���<T��<V��<j��<���<v��<���<���<��<���<`   `   *��<l��<[��<���<b��<r��<���<Z��<���<i��<���<���<���<���<���<i��<���<Z��<���<r��<b��<���<[��<l��<`   `   N��<���<p��<]��<k��<���<a��<F��<Ӟ�<���<���<���<c��<���<���<���<Ӟ�<F��<a��<���<k��<]��<p��<���<`   `   ���<���<}��<��<���<���<\��<w��<���<o��<���<}��<���<}��<���<o��<���<w��<\��<���<���<��<}��<���<`   `   ���<`��<���<���<w��<n��<���<ў�<y��<���<���<t��<���<t��<���<���<y��<ў�<���<n��<w��<���<���<`��<`   `   ў�<���<���<z��<@��<R��<s��<���<~��<���<��<b��<���<b��<��<���<~��<���<s��<R��<@��<z��<���<���<`   `   ���<���<���<���<���<_��<[��<���<���<���<��<���<���<���<��<���<���<���<[��<_��<���<���<���<���<`   `   z��<��<`��<���<���<���<���<���<���<��<���<���<e��<���<���<��<���<���<���<���<���<���<`��<��<`   `   ��<˞�<���<���<���<ɞ�<���<���<���<f��<���<}��<~��<}��<���<f��<���<���<���<ɞ�<���<���<���<˞�<`   `   ߞ�<���<���<۞�<���<���<���<���<���<���<���<t��<���<t��<���<���<���<���<���<���<���<۞�<���<���<`   `   ��<���<���<۞�<���<���<���<���<���<���<���<b��<y��<b��<���<���<���<���<���<���<���<۞�<���<���<`   `   Ξ�<Ǟ�<���<���<}��<j��<���<���<���<g��<���<���<k��<���<���<g��<���<���<���<j��<}��<���<���<Ǟ�<`   `   q��<���<Ӟ�<���<���<���<���<Þ�<���<X��<���<���<p��<���<���<X��<���<Þ�<���<���<���<���<Ӟ�<���<`   `   ɞ�<��<��<Þ�<Þ�<؞�<���<���<���<Q��<���<p��<G��<p��<���<Q��<���<���<���<؞�<Þ�<Þ�<��<��<`   `   	��<˞�<���<���<���<ٞ�<���<���<���<A��<n��<U��<y��<U��<n��<A��<���<���<���<ٞ�<���<���<���<˞�<`   `   מ�<���<���<���<���<���<d��<x��<y��<N��<���<���<���<���<���<N��<y��<x��<d��<���<���<���<���<���<`   `   ɞ�<���<���<���<Ǟ�<���<x��<���<���<v��<���<v��<]��<v��<���<v��<���<���<x��<���<Ǟ�<���<���<���<`   `   ��<Ş�<���<���<Ϟ�<���<���<˞�<���<|��<X��<]��<���<]��<X��<|��<���<˞�<���<���<Ϟ�<���<���<Ş�<`   `   ƞ�<���<���<���<���<��<���<���<k��<���<d��<z��<Ϟ�<z��<d��<���<k��<���<���<��<���<���<���<���<`   `   ���<���<Ξ�<���<���<���<Þ�<���<���<���<y��<N��<��<N��<y��<���<���<���<Þ�<���<���<���<Ξ�<���<`   `   n��<���<���<���<���<y��<���<n��<���<h��<7��<{��<H��<{��<7��<h��<���<n��<���<y��<���<���<���<���<`   `   K��<���<���<���<���<v��<���<z��<���<V��<Y��<���<^��<���<Y��<V��<���<z��<���<v��<���<���<���<���<`   `   ���<�<���<���<���<N��<���<���<z��<k��<���<l��<֝�<l��<���<k��<z��<���<���<N��<���<���<���<�<`   `   ���<���<���<���<=��<D��<���<z��<r��<Y��<*��<j��<I��<j��<*��<Y��<r��<z��<���<D��<=��<���<���<���<`   `   ���<~��<���<T��<V��<j��<���<v��<���<���<��<���<���<���<��<���<���<v��<���<j��<V��<T��<���<~��<`   `   ���<���<���<i��<���<Z��<���<r��<b��<���<[��<l��<*��<l��<[��<���<b��<r��<���<Z��<���<i��<���<���<`   `   c��<���<���<���<Ӟ�<F��<a��<���<k��<]��<p��<���<N��<���<p��<]��<k��<���<a��<F��<Ӟ�<���<���<���<`   `   ���<}��<���<o��<���<w��<\��<���<���<��<}��<���<���<���<}��<��<���<���<\��<w��<���<o��<���<}��<`   `   ���<t��<���<���<y��<ў�<���<n��<w��<���<���<`��<���<`��<���<���<w��<n��<���<ў�<y��<���<���<t��<`   `   ���<b��<��<���<}��<���<s��<R��<@��<z��<���<���<ў�<���<���<z��<@��<R��<s��<���<}��<���<��<b��<`   `   ���<���<��<���<���<���<[��<_��<���<���<���<���<���<���<���<���<���<_��<[��<���<���<���<��<���<`   `   e��<���<���<��<���<���<���<���<���<���<`��<��<z��<��<`��<���<���<���<���<���<���<��<���<���<`   `   ~��<}��<���<f��<���<���<���<ɞ�<���<���<���<˞�<��<˞�<���<���<���<ɞ�<���<���<���<f��<���<}��<`   `   ���<t��<���<���<���<���<���<���<���<۞�<���<���<ߞ�<���<���<۞�<���<���<���<���<���<���<���<t��<`   `   y��<b��<���<���<���<���<���<���<���<۞�<���<���<��<���<���<۞�<���<���<���<���<���<���<���<b��<`   `   k��<���<���<g��<���<���<���<j��<}��<���<���<Ǟ�<Ξ�<Ǟ�<���<���<}��<j��<���<���<���<g��<���<���<`   `   p��<���<���<X��<���<Þ�<���<���<���<���<Ӟ�<���<q��<���<Ӟ�<���<���<���<���<Þ�<���<X��<���<���<`   `   G��<p��<���<Q��<���<���<���<؞�<Þ�<Þ�<��<��<ɞ�<��<��<Þ�<Þ�<؞�<���<���<���<Q��<���<p��<`   `   y��<U��<n��<A��<���<���<���<ٞ�<���<���<���<˞�<	��<˞�<���<���<���<ٞ�<���<���<���<A��<n��<U��<`   `   ���<���<���<N��<y��<x��<d��<���<���<���<���<���<מ�<���<���<���<���<���<d��<x��<y��<N��<���<���<`   `   ]��<v��<���<v��<���<���<x��<���<Ǟ�<���<���<���<ɞ�<���<���<���<Ǟ�<���<x��<���<���<v��<���<v��<`   `   ���<]��<X��<|��<���<̞�<���<���<Ϟ�<���<���<Ş�<��<Ş�<���<���<Ϟ�<���<���<̞�<���<|��<X��<]��<`   `   Ϟ�<z��<d��<���<k��<���<���<��<���<���<���<���<ƞ�<���<���<���<���<��<���<���<k��<���<d��<z��<`   `   ��<N��<y��<���<���<���<Þ�<���<���<���<Ξ�<���<���<���<Ξ�<���<���<���<Þ�<���<���<���<y��<N��<`   `   H��<{��<7��<h��<���<n��<���<y��<���<���<���<���<n��<���<���<���<���<y��<���<n��<���<h��<7��<{��<`   `   ^��<���<Y��<V��<���<z��<���<v��<���<���<���<���<K��<���<���<���<���<v��<���<z��<���<V��<Y��<���<`   `   ��<|��<���<���<w��<~��<���<���<���<y��<���<Ѡ�<Ǡ�<Ѡ�<���<y��<���<���<���<~��<w��<���<���<|��<`   `   ���<���<���<j��<h��<q��<M��< �<��<���<���<���<���<���<���<���<��< �<M��<q��<h��<j��<���<���<`   `   ?��<���<���<o��<���<���<���<Ơ�<��<Ġ�<���<u��<à�<u��<���<Ġ�<��<Ơ�<���<���<���<o��<���<���<`   `   n��<���<t��<}��<d��<]��<���<���<h��<���<���<���<͠�<���<���<���<h��<���<���<]��<d��<}��<t��<���<`   `   <��<v��<Z��<���<���<c��<���<���<j��<v��<���<���<���<���<���<v��<j��<���<���<c��<���<���<Z��<v��<`   `   o��<���<���<���<���<���<���<Ѡ�<���<���<���<���<���<���<���<���<���<Ѡ�<���<���<���<���<���<���<`   `   ���<{��<���<p��<s��<���<J��<\��<���<���<���<���<���<���<���<���<���<\��<J��<���<s��<p��<���<{��<`   `   n��<I��<���<���<Π�<
��<���<j��<���<~��<���<���<���<���<���<~��<���<j��<���<
��<Π�<���<���<I��<`   `   Ϡ�<���<���<���<���<Р�<ܠ�<���<���<���<���<���<x��<���<���<���<���<���<ܠ�<Р�<���<���<���<���<`   `   ���<Ϡ�<���<���<|��<z��<���<z��<���<���<���<���<w��<���<���<���<���<z��<���<z��<|��<���<���<Ϡ�<`   `   p��<���<ɠ�<��<���<���<~��<|��<���<x��<���<���<���<���<���<x��<���<|��<~��<���<���<��<ɠ�<���<`   `   ̠�<���<Ӡ�<��<v��<���<���<���<���<���<���<v��<���<v��<���<���<���<���<���<���<v��<��<Ӡ�<���<`   `   ���<ڠ�<Ǡ�<��<���<Ԡ�<ʠ�<���<n��<���<̠�<v��<���<v��<̠�<���<n��<���<ʠ�<Ԡ�<���<��<Ǡ�<ڠ�<`   `   Ƞ�<Ӡ�<Ġ�<Ǡ�<��<��<Ǡ�<���<{��<���<���<���<Р�<���<���<���<{��<���<Ǡ�<��<��<Ǡ�<Ġ�<Ӡ�<`   `   ���<ݠ�<���<���<ܠ�<Ԡ�<m��<���<���<Ѡ�<t��<j��<ˠ�<j��<t��<Ѡ�<���<���<m��<Ԡ�<ܠ�<���<���<ݠ�<`   `   ޠ�<��<!��<���<���<Š�<~��<z��<���<��<���<}��<ڠ�<}��<���<��<���<z��<~��<Š�<���<���<!��<��<`   `   ��<ˠ�<��<��<Ϡ�<��<��<���<���<��<���<���<���<���<���<��<���<���<��<��<Ϡ�<��<��<ˠ�<`   `    ��<���<Ҡ�<���<Ƞ�<���<ڠ�<���<٠�<���<���<���<1��<���<���<���<٠�<���<ڠ�<���<Ƞ�<���<Ҡ�<���<`   `    ��<��<ߠ�<���<Ԡ�<���<���<���<Ԡ�<���<c��<���<'��<���<c��<���<Ԡ�<���<���<���<Ԡ�<���<ߠ�<��<`   `   ��<���<Ӡ�<Ӡ�<Ƞ�<���<Ҡ�<g��<���<���<��<���<b��<���<��<���<���<g��<Ҡ�<���<Ƞ�<Ӡ�<Ӡ�<���<`   `   ���<���<ɠ�<���<���<���<���<Q��<���<���<���<e��<V��<e��<���<���<���<Q��<���<���<���<���<ɠ�<���<`   `   ���<Ԡ�<ޠ�<��<���<ɠ�<|��<o��<���<m��<���<���<���<���<���<m��<���<o��<|��<ɠ�<���<��<ޠ�<Ԡ�<`   `   ��<Ҡ�<���<��<̠�< �<m��<���<|��<=��<���<���<���<���<���<=��<|��<���<m��< �<̠�<��<���<Ҡ�<`   `   Ǡ�<���<t��<���<���<Ġ�<���<���<���<���<���<G��<���<G��<���<���<���<���<���<Ġ�<���<���<t��<���<`   `   Ǡ�<Ѡ�<���<y��<���<���<���<~��<w��<���<���<|��<��<|��<���<���<w��<~��<���<���<���<y��<���<Ѡ�<`   `   ���<���<���<���<��< �<M��<q��<h��<j��<���<���<���<���<���<j��<h��<q��<M��< �<��<���<���<���<`   `   à�<u��<���<Ġ�<��<Ơ�<���<���<���<o��<���<���<?��<���<���<o��<���<���<���<Ơ�<��<Ġ�<���<u��<`   `   ͠�<���<���<���<h��<���<���<]��<d��<}��<t��<���<n��<���<t��<}��<d��<]��<���<���<h��<���<���<���<`   `   ���<���<���<v��<j��<���<���<c��<���<���<Z��<v��<<��<v��<Z��<���<���<c��<���<���<j��<v��<���<���<`   `   ���<���<���<���<���<Ѡ�<���<���<���<���<���<���<o��<���<���<���<���<���<���<Ѡ�<���<���<���<���<`   `   ���<���<���<���<���<\��<J��<���<s��<p��<���<{��<���<{��<���<p��<s��<���<J��<\��<���<���<���<���<`   `   ���<���<���<~��<���<j��<���<
��<Π�<���<���<I��<n��<I��<���<���<Π�<
��<���<j��<���<~��<���<���<`   `   x��<���<���<���<���<���<ܠ�<Р�<���<���<���<���<Ϡ�<���<���<���<���<Р�<ܠ�<���<���<���<���<���<`   `   w��<���<���<���<���<z��<���<z��<|��<���<���<Ϡ�<���<Ϡ�<���<���<|��<z��<���<z��<���<���<���<���<`   `   ���<���<���<x��<���<|��<~��<���<���<��<ɠ�<���<p��<���<ɠ�<��<���<���<~��<|��<���<x��<���<���<`   `   ���<v��<���<���<���<���<���<���<v��<��<Ӡ�<���<̠�<���<Ӡ�<��<v��<���<���<���<���<���<���<v��<`   `   ���<v��<̠�<���<n��<���<ʠ�<Ԡ�<���<��<Ǡ�<ڠ�<���<ڠ�<Ǡ�<��<���<Ԡ�<ʠ�<���<n��<���<̠�<v��<`   `   Р�<���<���<���<{��<���<Ǡ�<��<��<Ǡ�<Ġ�<Ӡ�<Ƞ�<Ӡ�<Ġ�<Ǡ�<��<��<Ǡ�<���<{��<���<���<���<`   `   ˠ�<j��<t��<Ѡ�<���<���<m��<Ԡ�<ܠ�<���<���<ݠ�<���<ݠ�<���<���<ܠ�<Ԡ�<m��<���<���<Ѡ�<t��<j��<`   `   ڠ�<}��<���<��<���<z��<~��<Š�<���<���<!��<��<ޠ�<��<!��<���<���<Š�<~��<z��<���<��<���<}��<`   `   ���<���<���<��<���<���<��<��<Ϡ�<��<��<ˠ�<��<ˠ�<��<��<Ϡ�<��<��<���<���<��<���<���<`   `   1��<���<���<���<٠�<���<ڠ�<���<Ƞ�<���<Ҡ�<���< ��<���<Ҡ�<���<Ƞ�<���<ڠ�<���<٠�<���<���<���<`   `   '��<���<c��<���<Ԡ�<���<���<���<Ԡ�<���<ߠ�<��< ��<��<ߠ�<���<Ԡ�<���<���<���<Ԡ�<���<c��<���<`   `   b��<���<��<���<���<g��<Ҡ�<���<Ƞ�<Ӡ�<Ӡ�<���<��<���<Ӡ�<Ӡ�<Ƞ�<���<Ҡ�<g��<���<���<��<���<`   `   V��<e��<���<���<���<Q��<���<���<���<���<ɠ�<���<���<���<ɠ�<���<���<���<���<Q��<���<���<���<e��<`   `   ���<���<���<m��<���<o��<|��<ɠ�<���<��<ޠ�<Ԡ�<���<Ԡ�<ޠ�<��<���<ɠ�<|��<o��<���<m��<���<���<`   `   ���<���<���<=��<|��<���<m��< �<̠�<��<���<Ҡ�<��<Ҡ�<���<��<̠�< �<m��<���<|��<=��<���<���<`   `   ���<G��<���<���<���<���<���<Ġ�<���<���<t��<���<Ǡ�<���<t��<���<���<Ġ�<���<���<���<���<���<G��<`   `   ��<K��<Q��<���<���<���<���<��<���<��<
��<��<Ģ�<��<
��<��<���<��<���<���<���<���<Q��<K��<`   `   k��<X��<���<���<���<Ģ�<���<���<���<���<��<��<���<��<��<���<���<���<���<Ģ�<���<���<���<X��<`   `   ��<T��<���<���<���<Ӣ�<~��<���<���<���<��<��<ߢ�<��<��<���<���<���<~��<Ӣ�<���<���<���<T��<`   `   ���<���<���<���<���<���<���<���<���<��<���<���<ˢ�<���<���<��<���<���<���<���<���<���<���<���<`   `   â�<���<���<ɢ�<Ǣ�<���<���<���<���<ޢ�<���<���<��<���<���<ޢ�<���<���<���<���<Ǣ�<ɢ�<���<���<`   `   ���<��<���<���<���<���<Ǣ�<���<���<Ģ�<���<Ţ�<٢�<Ţ�<���<Ģ�<���<���<Ǣ�<���<���<���<���<��<`   `   %��<��<���<���<���<���<¢�<���<���<���<���<���<|��<���<���<���<���<���<¢�<���<���<���<���<��<`   `   ݢ�<̢�<���<Ң�<Ǣ�<{��<���<آ�<֢�<ˢ�<���<̢�<���<̢�<���<ˢ�<֢�<آ�<���<{��<Ǣ�<Ң�<���<̢�<`   `   ���<٢�<Ƣ�<���<���<~��<ʢ�<Ǣ�<���<Ϣ�<���<���<ɢ�<���<���<Ϣ�<���<Ǣ�<ʢ�<~��<���<���<Ƣ�<٢�<`   `   ߢ�<	��<��<���<��<ɢ�<��<Ţ�<���<��<���<���<¢�<���<���<��<���<Ţ�<��<ɢ�<��<���<��<	��<`   `   ��<��<ۢ�<Ԣ�<9��< ��<���<��<���<��<֢�<���<���<���<֢�<��<���<��<���< ��<9��<Ԣ�<ۢ�<��<`   `   ���<.��<��<���<��<��<Ȣ�<ߢ�<͢�<���<���<���<���<���<���<���<͢�<ߢ�<Ȣ�<��<��<���<��<.��<`   `   ���<��<��<ݢ�<��<ע�<���<Ǣ�<��<���<���<���<Ң�<���<���<���<��<Ǣ�<���<ע�<��<ݢ�<��<��<`   `   #��<&��</��<0��<��<Ȣ�<��<��<��<Ȣ�<���<���<���<���<���<Ȣ�<��<��<��<Ȣ�<��<0��</��<&��<`   `   ���<=��<���<,��<���<��<6��<��<���<���<���<���<u��<���<���<���<���<��<6��<��<���<,��<���<=��<`   `   ?��<Т�<͢�<��<��<Ң�<��<'��<���<���<���<΢�<���<΢�<���<���<���<'��<��<Ң�<��<��<͢�<Т�<`   `   ��<	��<8��<$��<1��<���<ˢ�<��<���<���<���<â�<���<â�<���<���<���<��<ˢ�<���<1��<$��<8��<	��<`   `   	��<b��<d��<բ�<'��<��<��<���<���<���<c��<���<���<���<c��<���<���<���<��<��<'��<բ�<d��<b��<`   `   Ǣ�<.��<��<���<���<��<��<â�<���<���<q��<��<΢�<��<q��<���<���<â�<��<��<���<���<��<.��<`   `   ߢ�< ��<��<��<��<��<��<Ң�<���<���<���<Ң�<���<Ң�<���<���<���<Ң�<��<��<��<��<��< ��<`   `   ��<+��<$��<#��<!��<��<���<��<ۢ�<v��<���<���<t��<���<���<v��<ۢ�<��<���<��<!��<#��<$��<+��<`   `   ��<��<͢�<���<��<��<â�<��<��<\��<}��<���<��<���<}��<\��<��<��<â�<��<��<���<͢�<��<`   `   ڢ�<��<٢�<բ�<���<Ѣ�<���<Ӣ�<���<���<��<_��<���<_��<��<���<���<Ӣ�<���<Ѣ�<���<բ�<٢�<��<`   `   բ�<��<(��<2��<���<���<���<���<m��<���<���<��<h��<��<���<���<m��<���<���<���<���<2��<(��<��<`   `   Ģ�<��<
��<��<���<��<���<���<���<���<Q��<K��<��<K��<Q��<���<���<���<���<��<���<��<
��<��<`   `   ���<��<��<���<���<���<���<Ģ�<���<���<���<X��<k��<X��<���<���<���<Ģ�<���<���<���<���<��<��<`   `   ߢ�<��<��<���<���<���<~��<Ӣ�<���<���<���<T��<��<T��<���<���<���<Ӣ�<~��<���<���<���<��<��<`   `   ˢ�<���<���<��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<��<���<���<`   `   ��<���<���<ޢ�<���<���<���<���<Ǣ�<ɢ�<���<���<â�<���<���<ɢ�<Ǣ�<���<���<���<���<ޢ�<���<���<`   `   ٢�<Ţ�<���<Ģ�<���<���<Ǣ�<���<���<���<���<��<���<��<���<���<���<���<Ǣ�<���<���<Ģ�<���<Ţ�<`   `   |��<���<���<���<���<���<¢�<���<���<���<���<��<%��<��<���<���<���<���<¢�<���<���<���<���<���<`   `   ���<̢�<���<ˢ�<֢�<آ�<���<{��<Ǣ�<Ң�<���<̢�<ݢ�<̢�<���<Ң�<Ǣ�<{��<���<آ�<֢�<ˢ�<���<̢�<`   `   ɢ�<���<���<Ϣ�<���<Ǣ�<ʢ�<~��<���<���<Ƣ�<٢�<���<٢�<Ƣ�<���<���<~��<ʢ�<Ǣ�<���<Ϣ�<���<���<`   `   ¢�<���<���<��<���<Ţ�<��<ɢ�<��<���<��<	��<ߢ�<	��<��<���<��<ɢ�<��<Ţ�<���<��<���<���<`   `   ���<���<֢�<��<���<��<���< ��<9��<Ԣ�<ۢ�<��<��<��<ۢ�<Ԣ�<9��< ��<���<��<���<��<֢�<���<`   `   ���<���<���<���<͢�<ߢ�<Ȣ�<��<��<���<��<.��<���<.��<��<���<��<��<Ȣ�<ߢ�<͢�<���<���<���<`   `   Ң�<���<���<���<��<Ǣ�<���<ע�<��<ݢ�<��<��<���<��<��<ݢ�<��<ע�<���<Ǣ�<��<���<���<���<`   `   ���<���<���<Ȣ�<��<��<��<Ȣ�<��<0��</��<&��<#��<&��</��<0��<��<Ȣ�<��<��<��<Ȣ�<���<���<`   `   u��<���<���<���<���<��<6��<��<���<,��<���<=��<���<=��<���<,��<���<��<6��<��<���<���<���<���<`   `   ���<΢�<���<���<���<'��<��<Ң�<��<��<͢�<Т�<?��<Т�<͢�<��<��<Ң�<��<'��<���<���<���<΢�<`   `   ���<â�<���<���<���<��<ˢ�<���<1��<$��<8��<	��<��<	��<8��<$��<1��<���<ˢ�<��<���<���<���<â�<`   `   ���<���<c��<���<���<���<��<��<'��<բ�<d��<b��<	��<b��<d��<բ�<'��<��<��<���<���<���<c��<���<`   `   ΢�<��<q��<���<���<â�<��<��<���<���<��<.��<Ǣ�<.��<��<���<���<��<��<â�<���<���<q��<��<`   `   ���<Ң�<���<���<���<Ң�<��<��<��<��<��< ��<ߢ�< ��<��<��<��<��<��<Ң�<���<���<���<Ң�<`   `   t��<���<���<v��<ۢ�<��<���<��<!��<#��<$��<+��<��<+��<$��<#��<!��<��<���<��<ۢ�<v��<���<���<`   `   ��<���<}��<\��<��<��<â�<��<��<���<͢�<��<��<��<͢�<���<��<��<â�<��<��<\��<}��<���<`   `   ���<_��<��<���<���<Ӣ�<���<Ѣ�<���<բ�<٢�<��<ڢ�<��<٢�<բ�<���<Ѣ�<���<Ӣ�<���<���<��<_��<`   `   h��<��<���<���<m��<���<���<���<���<2��<(��<��<բ�<��<(��<2��<���<���<���<���<m��<���<���<��<`   `   g��<ۤ�<���<{��<��<ɤ�<��<��<��<��<���<���<K��<���<���<��<��<��<��<ɤ�<��<{��<���<ۤ�<`   `   Ȥ�<ɤ�<���<���<���<���<��<��<���<��<��<��<��<��<��<��<���<��<��<���<���<���<���<ɤ�<`   `   ��<���<���<���<���<���<��<��<ܤ�<��<��<��<Ҥ�<��<��<��<ܤ�<��<��<���<���<���<���<���<`   `   ���<c��<���<���<���<Ӥ�<֤�<��<��<֤�<���<���<Ƥ�<���<���<֤�<��<��<֤�<Ӥ�<���<���<���<c��<`   `   ���<���<��<���<���<֤�<���<Ϥ�<��<��<��<��<��<��<��<��<��<Ϥ�<���<֤�<���<���<��<���<`   `   ���<���<��<���<֤�<��<���<���<��<ܤ�<ޤ�<���<���<���<ޤ�<ܤ�<��<���<���<��<֤�<���<��<���<`   `   ���<���<���<���<&��<���<��<��<��<ͤ�<Ƥ�<ߤ�<ɤ�<ߤ�<Ƥ�<ͤ�<��<��<��<���<&��<���<���<���<`   `   Ť�<���<��<��<���<Ĥ�<��<��<Ԥ�<٤�<��<��<��<��<��<٤�<Ԥ�<��<��<Ĥ�<���<��<��<���<`   `   ��<��<��<��<��<��<Ԥ�<Ȥ�<Ϥ�<��<ޤ�<פ�<��<פ�<ޤ�<��<Ϥ�<Ȥ�<Ԥ�<��<��<��<��<��<`   `   ��<ߤ�<��<%��<��<��<��<��<���<���<ͤ�<��<��<��<ͤ�<���<���<��<��<��<��<%��<��<ߤ�<`   `   >��<��<&��<5��<ڤ�<���<��<��<פ�<��<ݤ�<��<ݤ�<��<ݤ�<��<פ�<��<��<���<ڤ�<5��<&��<��<`   `   c��<H��<L��<U��<6��<��<��<��<ɤ�<���<��<���<���<���<��<���<ɤ�<��<��<��<6��<U��<L��<H��<`   `   c��<d��<C��<[��<s��<O��<R��<��<.��<��<ܤ�<��<���<��<ܤ�<��<.��<��<R��<O��<s��<[��<C��<d��<`   `   6��<<��<-��<B��<��<��<%��<��<��<��<ؤ�<���<���<���<ؤ�<��<��<��<%��<��<��<B��<-��<<��<`   `   '��<M��<o��<m��<3��<C��<��<���<��<��<	��<��<Ԥ�<��<	��<��<��<���<��<C��<3��<m��<o��<M��<`   `   a��<���<���<U��<V��<w��<��<��<6��<��<��<��<���<��<��<��<6��<��<��<w��<V��<U��<���<���<`   `   ���<���<m��<��<6��<F��<��<��<!��<��<ޤ�<դ�<���<դ�<ޤ�<��<!��<��<��<F��<6��<��<m��<���<`   `   ���<J��<N��<V��<q��<A��<��< ��<��<$��<��<��<դ�<��<��<$��<��< ��<��<A��<q��<V��<N��<J��<`   `   ���<:��<k��<���<r��<��<��<��<ڤ�<��<ؤ�<���<���<���<ؤ�<��<ڤ�<��<��<��<r��<���<k��<:��<`   `   ���<;��<M��<{��<'��<���<��<��<Ӥ�<Ϥ�<¤�<y��<���<y��<¤�<Ϥ�<Ӥ�<��<��<���<'��<{��<M��<;��<`   `   {��<:��<(��<J��<��<��<��<Ҥ�<���<��<���<���<Ǥ�<���<���<��<���<Ҥ�<��<��<��<J��<(��<:��<`   `   
��<W��<V��<A��<��<��<��<���<���<��<���<v��<���<v��<���<��<���<���<��<��<��<A��<V��<W��<`   `   ��<Z��<Q��<��<,��<��<��<ä�<Ĥ�<Ȥ�<���<���<���<���<���<Ȥ�<Ĥ�<ä�<��<��<,��<��<Q��<Z��<`   `   P��<7��<��<���<��<��<ݤ�<Ǥ�<٤�<���<Ƥ�<��<���<��<Ƥ�<���<٤�<Ǥ�<ݤ�<��<��<���<��<7��<`   `   K��<���<���<��<��<��<��<ɤ�<��<{��<���<ۤ�<g��<ۤ�<���<{��<��<ɤ�<��<��<��<��<���<���<`   `   ��<��<��<��<���<��<��<���<���<���<���<ɤ�<Ȥ�<ɤ�<���<���<���<���<��<��<���<��<��<��<`   `   Ҥ�<��<��<��<ܤ�<��<��<���<���<���<���<���<��<���<���<���<���<���<��<��<ܤ�<��<��<��<`   `   Ƥ�<���<���<֤�<��<��<֤�<Ӥ�<���<���<���<c��<���<c��<���<���<���<Ӥ�<֤�<��<��<֤�<���<���<`   `   ��<��<��<��<��<Ϥ�<���<֤�<���<���<��<���<���<���<��<���<���<֤�<���<Ϥ�<��<��<��<��<`   `   ���<���<ޤ�<ܤ�<��<���<���<��<֤�<���<��<���<���<���<��<���<֤�<��<���<���<��<ܤ�<ޤ�<���<`   `   ɤ�<ߤ�<Ƥ�<ͤ�<��<��<��<���<&��<���<���<���<���<���<���<���<&��<���<��<��<��<ͤ�<Ƥ�<ߤ�<`   `   ��<��<��<٤�<Ԥ�<��<��<Ĥ�<���<��<��<���<Ť�<���<��<��<���<Ĥ�<��<��<Ԥ�<٤�<��<��<`   `   ��<פ�<ޤ�<��<Ϥ�<Ȥ�<Ԥ�<��<��<��<��<��<��<��<��<��<��<��<Ԥ�<Ȥ�<Ϥ�<��<ޤ�<פ�<`   `   ��<��<ͤ�<���<���<��<��<��<��<%��<��<ߤ�<��<ߤ�<��<%��<��<��<��<��<���<���<ͤ�<��<`   `   ݤ�<��<ݤ�<��<פ�<��<��<���<ڤ�<5��<&��<��<>��<��<&��<5��<ڤ�<���<��<��<פ�<��<ݤ�<��<`   `   ���<���<��<���<ɤ�<��<��<��<6��<U��<L��<H��<c��<H��<L��<U��<6��<��<��<��<ɤ�<���<��<���<`   `   ���<��<ܤ�<��<.��<��<R��<O��<s��<[��<C��<d��<c��<d��<C��<[��<s��<O��<R��<��<.��<��<ܤ�<��<`   `   ���<���<ؤ�<��<��<��<%��<��<��<B��<-��<<��<6��<<��<-��<B��<��<��<%��<��<��<��<ؤ�<���<`   `   Ԥ�<��<	��<��<��<���<��<C��<3��<m��<o��<M��<'��<M��<o��<m��<3��<C��<��<���<��<��<	��<��<`   `   ���<��<��<��<6��<��<��<w��<V��<U��<���<���<a��<���<���<U��<V��<w��<��<��<6��<��<��<��<`   `   ���<դ�<ޤ�<��<!��<��<��<F��<6��<��<m��<���<���<���<m��<��<6��<F��<��<��<!��<��<ޤ�<դ�<`   `   դ�<��<��<$��<��< ��<��<A��<q��<V��<N��<J��<���<J��<N��<V��<q��<A��<��< ��<��<$��<��<��<`   `   ���<���<ؤ�<��<ڤ�<��<��<��<r��<���<k��<:��<���<:��<k��<���<r��<��<��<��<ڤ�<��<ؤ�<���<`   `   ���<y��<¤�<Ϥ�<Ӥ�<��<��<���<'��<{��<M��<;��<���<;��<M��<{��<'��<���<��<��<Ӥ�<Ϥ�<¤�<y��<`   `   Ǥ�<���<���<��<���<Ҥ�<��<��<��<J��<(��<:��<{��<:��<(��<J��<��<��<��<Ҥ�<���<��<���<���<`   `   ���<v��<���<��<���<���<��<��<��<A��<V��<W��<
��<W��<V��<A��<��<��<��<���<���<��<���<v��<`   `   ���<���<���<Ȥ�<Ĥ�<ä�<��<��<,��<��<Q��<Z��<��<Z��<Q��<��<,��<��<��<ä�<Ĥ�<Ȥ�<���<���<`   `   ���<��<Ƥ�<���<٤�<Ǥ�<ݤ�<��<��<���<��<7��<P��<7��<��<���<��<��<ݤ�<Ǥ�<٤�<���<Ƥ�<��<`   `   ��<���<���<��<��<˦�<��<��<'��<@��<���<m��<Y��<m��<���<@��<'��<��<��<˦�<��<��<���<���<`   `   ��<���<���<��<��<��<��<��<@��<X��<P��<Z��<C��<Z��<P��<X��<@��<��<��<��<��<��<���<���<`   `   ��<��<Ʀ�<��<��<צ�<���<��<+��<J��<��<@��<)��<@��<��<J��<+��<��<���<צ�<��<��<Ʀ�<��<`   `   x��<���<��<���<��<���<���<��<Ӧ�<#��<4��<N��<��<N��<4��<#��<Ӧ�<��<���<���<��<���<��<���<`   `   ��<��<���<���<ۦ�<��<��<��<ͦ�<���<5��<6��<��<6��<5��<���<ͦ�<��<��<��<ۦ�<���<���<��<`   `   F��<��<ݦ�<��<��<��<��<*��<&��<��<��<��<��<��<��<��<&��<*��<��<��<��<��<ݦ�<��<`   `   ���<��<���<��<��<��<��<ަ�<��</��<��<#��<h��<#��<��</��<��<ަ�<��<��<��<��<���<��<`   `   ,��<P��<,��<��<��<+��<"��<���<��<��<��<���<,��<���<��<��<��<���<"��<+��<��<��<,��<P��<`   `   ���<;��<C��<>��<��<y��<6��<@��<J��<��<<��<���<���<���<<��<��<J��<@��<6��<y��<��<>��<C��<;��<`   `   ӧ�<]��<z��<]��</��<���<��<*��<G��<���<9��<D��<��<D��<9��<���<G��<*��<��<���</��<]��<z��<]��<`   `   ���<o��<���<`��<O��<���<\��<0��<?��<��<��<��<��<��<��<��<?��<0��<\��<���<O��<`��<���<o��<`   `   c��<Y��<���<|��<u��<t��<}��<4��<4��<N��<���<+��<��<+��<���<N��<4��<4��<}��<t��<u��<|��<���<Y��<`   `   ��<���<���<���<���<g��<l��<D��<��<0��<��<%��<��<%��<��<0��<��<D��<l��<g��<���<���<���<���<`   `   ��<���<���<���<���<���<y��<���<'��<��<
��<��<��<��<
��<��<'��<���<y��<���<���<���<���<���<`   `   ���<��<§�<���<���<���<p��<���<X��<A��<��<Ц�<Q��<Ц�<��<A��<X��<���<p��<���<���<���<§�<��<`   `   ���<���<֧�<���<���<���<`��<>��<[��<D��<��<��<D��<��<��<D��<[��<>��<`��<���<���<���<֧�<���<`   `   ̧�<ȧ�<ħ�<��<��<���<���<(��<'��<���<���< ��<2��< ��<���<���<'��<(��<���<���<��<��<ħ�<ȧ�<`   `   ��<���<���<��<f��<���<���<t��<��<ئ�<���<��<��<��<���<ئ�<��<t��<���<���<f��<��<���<���<`   `   ��<ק�<��<���<A��<{��<7��<N��<��<��<���<ܦ�<)��<ܦ�<���<��<��<N��<7��<{��<A��<���<��<ק�<`   `   ŧ�<���<ϧ�<q��<[��<��<b��<5��<0��<Φ�<Φ�<��<1��<��<Φ�<Φ�<0��<5��<b��<��<[��<q��<ϧ�<���<`   `   ���<���<���<p��<x��<ħ�<���<9��<-��<��<ߦ�<��<��<��<ߦ�<��<-��<9��<���<ħ�<x��<p��<���<���<`   `   ���<���<���<���<���<��<N��<��<��<
��<ܦ�<��<���<��<ܦ�<
��<��<��<N��<��<���<���<���<���<`   `   ���<���<j��<b��<���<)��<M��<��<��<Ѧ�<y��<֦�<���<֦�<y��<Ѧ�<��<��<M��<)��<���<b��<j��<���<`   `   w��<s��<v��<��<J��<9��<��<��<��<¦�<���<���<x��<���<���<¦�<��<��<��<9��<J��<��<v��<s��<`   `   Y��<m��<���<@��<'��<��<��<˦�<��<��<���<���<��<���<���<��<��<˦�<��<��<'��<@��<���<m��<`   `   C��<Z��<P��<X��<@��<��<��<��<��<��<���<���<��<���<���<��<��<��<��<��<@��<X��<P��<Z��<`   `   )��<@��<��<J��<+��<��<���<צ�<��<��<Ʀ�<��<��<��<Ʀ�<��<��<צ�<���<��<+��<J��<��<@��<`   `   ��<N��<4��<#��<Ӧ�<��<���<���<��<���<��<���<x��<���<��<���<��<���<���<��<Ӧ�<#��<4��<N��<`   `   ��<6��<5��<���<ͦ�<��<��<��<ۦ�<���<���<��<��<��<���<���<ۦ�<��<��<��<ͦ�<���<5��<6��<`   `   ��<��<��<��<&��<*��<��<��<��<��<ݦ�<��<F��<��<ݦ�<��<��<��<��<*��<&��<��<��<��<`   `   h��<#��<��</��<��<ަ�<��<��<��<��<���<��<���<��<���<��<��<��<��<ަ�<��</��<��<#��<`   `   ,��<���<��<��<��<���<"��<+��<��<��<,��<P��<,��<P��<,��<��<��<+��<"��<���<��<��<��<���<`   `   ���<���<<��<��<J��<@��<6��<y��<��<>��<C��<;��<���<;��<C��<>��<��<y��<6��<@��<J��<��<<��<���<`   `   ��<D��<9��<���<G��<*��<��<���</��<]��<z��<]��<ӧ�<]��<z��<]��</��<���<��<*��<G��<���<9��<D��<`   `   ��<��<��<��<?��<0��<\��<���<O��<`��<���<o��<���<o��<���<`��<O��<���<\��<0��<?��<��<��<��<`   `   ��<+��<���<N��<4��<4��<}��<t��<u��<|��<���<Y��<c��<Y��<���<|��<u��<t��<}��<4��<4��<N��<���<+��<`   `   ��<%��<��<0��<��<D��<l��<g��<���<���<���<���<��<���<���<���<���<g��<l��<D��<��<0��<��<%��<`   `   ��<��<
��<��<'��<���<y��<���<���<���<���<���<��<���<���<���<���<���<y��<���<'��<��<
��<��<`   `   Q��<Ц�<��<A��<X��<���<p��<���<���<���<§�<��<���<��<§�<���<���<���<p��<���<X��<A��<��<Ц�<`   `   D��<��<��<D��<[��<>��<`��<���<���<���<֧�<���<���<���<֧�<���<���<���<`��<>��<[��<D��<��<��<`   `   2��< ��<���<���<'��<(��<���<���<��<��<ħ�<ȧ�<̧�<ȧ�<ħ�<��<��<���<���<(��<'��<���<���< ��<`   `   ��<��<���<ئ�<��<t��<���<���<f��<��<���<���<��<���<���<��<f��<���<���<t��<��<ئ�<���<��<`   `   )��<ܦ�<���<��<��<N��<7��<{��<A��<���<��<ק�<��<ק�<��<���<A��<{��<7��<N��<��<��<���<ܦ�<`   `   1��<��<Φ�<Φ�<0��<5��<b��<��<[��<q��<ϧ�<���<ŧ�<���<ϧ�<q��<[��<��<b��<5��<0��<Φ�<Φ�<��<`   `   ��<��<ߦ�<��<-��<9��<���<ħ�<x��<p��<���<���<���<���<���<p��<x��<ħ�<���<9��<-��<��<ߦ�<��<`   `   ���<��<ܦ�<
��<��<��<N��<��<���<���<���<���<���<���<���<���<���<��<N��<��<��<
��<ܦ�<��<`   `   ���<֦�<y��<Ѧ�<��<��<M��<)��<���<b��<j��<���<���<���<j��<b��<���<)��<M��<��<��<Ѧ�<y��<֦�<`   `   x��<���<���<¦�<��<��<��<9��<J��<��<v��<s��<w��<s��<v��<��<J��<9��<��<��<��<¦�<���<���<`   `   ���<��<��<%��<¨�<Z��<b��<���<���<���<��<���<���<���<��<���<���<���<b��<Z��<¨�<%��<��<��<`   `   ��<��<ը�<ڨ�<��<o��<F��<a��<f��<��<���<���<���<���<���<��<f��<a��<F��<o��<��<ڨ�<ը�<��<`   `   ���<��<��<���<���<+��<&��<n��<q��<[��<h��<���<���<���<h��<[��<q��<n��<&��<+��<���<���<��<��<`   `   ���<��<	��<̨�<��<���<(��<h��<d��<���<k��<O��<���<O��<k��<���<d��<h��<(��<���<��<̨�<	��<��<`   `   A��<��<ڨ�</��<2��<��<<��<R��<P��<���<H��<N��<���<N��<H��<���<P��<R��<<��<��<2��</��<ڨ�<��<`   `   
��<��<��<���<R��<;��<T��<`��<[��<K��<N��<O��<}��<O��<N��<K��<[��<`��<T��<;��<R��<���<��<��<`   `   ��<f��<`��<`��<B��<_��<_��<L��<F��<H��<r��<?��<\��<?��<r��<H��<F��<L��<_��<_��<B��<`��<`��<f��<`   `   ^��<���<V��<���<}��<z��<{��<y��<i��<O��<K��<��<o��<��<K��<O��<i��<y��<{��<z��<}��<���<V��<���<`   `   W��<O��<c��<��<���<,��<_��<���<q��<J��<M��<L��<���<L��<M��<J��<q��<���<_��<,��<���<��<c��<O��<`   `   ~��<���<���<���<���<A��<[��<Z��<1��<X��<j��<U��<^��<U��<j��<X��<1��<Z��<[��<A��<���<���<���<���<`   `   ک�<��<٩�<���<��<��<���<���<q��<���<Y��<E��<>��<E��<Y��<���<q��<���<���<��<��<���<٩�<��<`   `   ��<'��<��<٩�<��<���<���<���<���<x��<H��<j��<n��<j��<H��<x��<���<���<���<���<��<٩�<��<'��<`   `   ��<��<5��<��<���<���<r��<���<���<\��<i��<M��<>��<M��<i��<\��<���<���<r��<���<���<��<5��<��<`   `   
��<��<^��<A��<��<��<���<���<��<���<���<T��<x��<T��<���<���<��<���<���<��<��<A��<^��<��<`   `   t��<V��<��<,��<��<Ω�<é�<��<M��<X��<���<2��<���<2��<���<X��<M��<��<é�<Ω�<��<,��<��<V��<`   `   ���<\��<��<B��<��<ǩ�<��<��<G��<H��<���<0��<8��<0��<���<H��<G��<��<��<ǩ�<��<B��<��<\��<`   `   W��<���<B��<y��<G��<��<���<y��<���<���<���<S��<4��<S��<���<���<���<y��<���<��<G��<y��<B��<���<`   `   I��<���<K��<��<+��<���<���<���<���<^��<+��< ��<��< ��<+��<^��<���<���<���<���<+��<��<K��<���<`   `   ��<k��<��<��<2��<���<���<���<n��<i��<��<.��<��<.��<��<i��<n��<���<���<���<2��<��<��<k��<`   `   ٩�<G��<6��<-��<'��<���<R��<H��<h��<b��<[��<��<ި�<��<[��<b��<h��<H��<R��<���<'��<-��<6��<G��<`   `   ��<X��<A��<"��<���<t��<J��<a��<n��<���<Ǩ�<è�<���<è�<Ǩ�<���<n��<a��<J��<t��<���<"��<A��<X��<`   `   &��<��<��<ҩ�<ȩ�<z��<i��<h��<'��<���<��<1��<ߨ�<1��<��<���<'��<h��<i��<z��<ȩ�<ҩ�<��<��<`   `   ��<���<ة�<���<���<}��<U��<O��<���<,��<��<��<ʨ�<��<��<,��<���<O��<U��<}��<���<���<ة�<���<`   `   ��<���<)��<ة�<���<���<W��<A��<ܨ�<;��<ը�<Ȩ�<��<Ȩ�<ը�<;��<ܨ�<A��<W��<���<���<ة�<)��<���<`   `   ���<���<��<���<���<���<b��<Z��<¨�<%��<��<��<���<��<��<%��<¨�<Z��<b��<���<���<���<��<���<`   `   ���<���<���<��<f��<a��<F��<o��<��<ڨ�<ը�<��<��<��<ը�<ڨ�<��<o��<F��<a��<f��<��<���<���<`   `   ���<���<h��<[��<q��<n��<&��<+��<���<���<��<��<���<��<��<���<���<+��<&��<n��<q��<[��<h��<���<`   `   ���<O��<k��<���<d��<h��<(��<���<��<̨�<	��<��<���<��<	��<̨�<��<���<(��<h��<d��<���<k��<O��<`   `   ���<N��<H��<���<P��<R��<<��<��<2��</��<ڨ�<��<A��<��<ڨ�</��<2��<��<<��<R��<P��<���<H��<N��<`   `   }��<O��<N��<K��<[��<`��<T��<;��<R��<���<��<��<
��<��<��<���<R��<;��<T��<`��<[��<K��<N��<O��<`   `   \��<?��<r��<H��<F��<L��<_��<_��<B��<`��<`��<f��<��<f��<`��<`��<B��<_��<_��<L��<F��<H��<r��<?��<`   `   o��<��<K��<O��<i��<y��<{��<z��<}��<���<V��<���<^��<���<V��<���<}��<z��<{��<y��<i��<O��<K��<��<`   `   ���<L��<M��<J��<q��<���<_��<+��<���<��<c��<O��<W��<O��<c��<��<���<+��<_��<���<q��<J��<M��<L��<`   `   ^��<U��<j��<X��<1��<Z��<[��<A��<���<���<���<���<~��<���<���<���<���<A��<[��<Z��<1��<X��<j��<U��<`   `   >��<E��<Y��<���<q��<���<���<��<��<���<٩�<��<ک�<��<٩�<���<��<��<���<���<q��<���<Y��<E��<`   `   n��<j��<H��<x��<���<���<���<���<��<٩�<��<'��<��<'��<��<٩�<��<���<���<���<���<x��<H��<j��<`   `   >��<M��<i��<\��<���<���<r��<���<���<��<5��<��<��<��<5��<��<���<���<r��<���<���<\��<i��<M��<`   `   x��<T��<���<���<��<���<���<��<��<A��<^��<��<
��<��<^��<A��<��<��<���<���<��<���<���<T��<`   `   ���<2��<���<X��<M��<��<é�<Ω�<��<,��<��<V��<t��<V��<��<,��<��<Ω�<é�<��<M��<X��<���<2��<`   `   8��<0��<���<H��<G��<��<��<ǩ�<��<B��<��<\��<���<\��<��<B��<��<ǩ�<��<��<G��<H��<���<0��<`   `   4��<S��<���<���<���<y��<���<��<G��<y��<B��<���<W��<���<B��<y��<G��<��<���<y��<���<���<���<S��<`   `   ��< ��<+��<^��<���<���<���<���<+��<��<K��<���<I��<���<K��<��<+��<���<���<���<���<^��<+��< ��<`   `   ��<.��<��<i��<n��<���<���<���<2��<��<��<k��<��<k��<��<��<2��<���<���<���<n��<i��<��<.��<`   `   ި�<��<[��<b��<h��<H��<R��<���<'��<-��<6��<G��<٩�<G��<6��<-��<'��<���<R��<H��<h��<b��<[��<��<`   `   ���<è�<Ǩ�<���<n��<a��<J��<t��<���<"��<A��<X��<��<X��<A��<"��<���<t��<J��<a��<n��<���<Ǩ�<è�<`   `   ߨ�<1��<��<���<'��<h��<i��<z��<ȩ�<ҩ�<��<��<&��<��<��<ҩ�<ȩ�<z��<i��<h��<'��<���<��<1��<`   `   ʨ�<��<��<,��<���<O��<U��<}��<���<���<ة�<���<��<���<ة�<���<���<}��<U��<O��<���<,��<��<��<`   `   ��<Ȩ�<ը�<;��<ܨ�<A��<W��<���<���<ة�<)��<���<��<���<)��<ة�<���<���<W��<A��<ܨ�<;��<ը�<Ȩ�<`   `   ݪ�<Ū�<���<��<6��<|��<Y��<���<���<���<���<��<���<��<���<���<���<���<Y��<|��<6��<��<���<Ū�<`   `   ���<Ϊ�<"��<U��<>��<9��<+��<���<��<��< ��< ��<��< ��< ��<��<��<���<+��<9��<>��<U��<"��<Ϊ�<`   `   Ϊ�<��<,��<`��<^��<M��<j��<���<���<ū�<��<��<���<��<��<ū�<���<���<j��<M��<^��<`��<,��<��<`   `   +��<'��<%��<F��<\��<v��<���<���<w��<v��<���<���<���<���<���<v��<w��<���<���<v��<\��<F��<%��<'��<`   `   ?��<?��<N��<Q��<H��<}��<T��<J��<���<���<���<«�<ī�<«�<���<���<���<J��<T��<}��<H��<Q��<N��<?��<`   `   L��<x��<���<K��<8��<���<h��<]��<���<���<���<���<���<���<���<���<���<]��<h��<���<8��<K��<���<x��<`   `   r��<���<���<D��<c��<���<���<���<���<p��<ë�<���<`��<���<ë�<p��<���<���<���<���<c��<D��<���<���<`   `   ���<ͫ�<���<���<ɫ�<���<y��<���<���<���<���<���<���<���<���<���<���<���<y��<���<ɫ�<���<���<ͫ�<`   `   6��<R��<���<��<���< ��<��<���<���<«�<���<���<ƫ�<���<���<«�<���<���<��< ��<���<��<���<R��<`   `   ��<t��<@��<
��< ��<��<I��<��<���<ӫ�<���<o��<���<o��<���<ӫ�<���<��<I��<��< ��<
��<@��<t��<`   `   ��<@��<4��<=��<$��<���<���<��<���<«�<���<���<���<���<���<«�<���<��<���<���<$��<=��<4��<@��<`   `   ���<���<l��<���<M��<��<
��<��<���<���<ɫ�<«�<���<«�<ɫ�<���<���<��<
��<��<M��<���<l��<���<`   `   ��<���<���<���<m��<���<���<��<��<���<���<���<^��<���<���<���<��<��<���<���<m��<���<���<���<`   `   ��<���<���<���<n��<Ϭ�<U��<��<*��<Ы�<���<���<���<���<���<Ы�<*��<��<U��<Ϭ�<n��<���<���<���<`   `   ���<	��<��<Ĭ�<|��<{��<���<���<��<ȫ�<���<���<���<���<���<ȫ�<��<���<���<{��<|��<Ĭ�<��<	��<`   `   ��<��<��<ݬ�<���<���<f��<��<	��<���<w��<���<H��<���<w��<���<	��<��<f��<���<���<ݬ�<��<��<`   `   ʬ�<��<���<���<���<|��<G��<��<
��<���<���<���<���<���<���<���<
��<��<G��<|��<���<���<���<��<`   `   Ȭ�<��<��<���<���<>��<!��<��<ҫ�<���<K��<���<���<���<K��<���<ҫ�<��<!��<>��<���<���<��<��<`   `   ���<���<���<��<���<>��<���< ��<~��<X��<0��<M��<`��<M��<0��<X��<~��< ��<���<>��<���<��<���<���<`   `   ;��<��<��<Ĭ�<]��<��<x��<���<o��<}��<S��<K��<g��<K��<S��<}��<o��<���<x��<��<]��<Ĭ�<��<��<`   `   ۬�<���<w��<g��<3��<3��<8��<���<���<���<G��<8��<t��<8��<G��<���<���<���<8��<3��<3��<g��<w��<���<`   `   d��<���<���<K��<N��<���<��<���<c��<Q��<,��<��<_��<��<,��<Q��<c��<���<��<���<N��<K��<���<���<`   `   ���<��<���<C��<	��<��<���<���<[��<1��<��<Ҫ�<���<Ҫ�<��<1��<[��<���<���<��<	��<C��<���<��<`   `   ߬�<;��<
��<��<ث�<���<l��<���<\��<��<���<���<Ǫ�<���<���<��<\��<���<l��<���<ث�<��<
��<;��<`   `   ���<��<���<���<���<���<Y��<|��<6��<��<���<Ū�<ݪ�<Ū�<���<��<6��<|��<Y��<���<���<���<���<��<`   `   ��< ��< ��<��<��<���<+��<9��<>��<U��<"��<Ϊ�<���<Ϊ�<"��<U��<>��<9��<+��<���<��<��< ��< ��<`   `   ���<��<��<ū�<���<���<j��<M��<^��<`��<,��<��<Ϊ�<��<,��<`��<^��<M��<j��<���<���<ū�<��<��<`   `   ���<���<���<v��<w��<���<���<v��<\��<F��<%��<'��<+��<'��<%��<F��<\��<v��<���<���<w��<v��<���<���<`   `   ī�<«�<���<���<���<J��<T��<}��<H��<Q��<N��<?��<?��<?��<N��<Q��<H��<}��<T��<J��<���<���<���<«�<`   `   ���<���<���<���<���<]��<h��<���<8��<K��<���<x��<L��<x��<���<K��<8��<���<h��<]��<���<���<���<���<`   `   `��<���<ë�<p��<���<���<���<���<c��<D��<���<���<r��<���<���<D��<c��<���<���<���<���<p��<ë�<���<`   `   ���<���<���<���<���<���<y��<���<ɫ�<���<���<ͫ�<���<ͫ�<���<���<ɫ�<���<y��<���<���<���<���<���<`   `   ƫ�<���<���<«�<���<���<��< ��<���<��<���<R��<6��<R��<���<��<���< ��<��<���<���<«�<���<���<`   `   ���<o��<���<ӫ�<���<��<I��<��< ��<
��<@��<t��<��<t��<@��<
��< ��<��<I��<��<���<ӫ�<���<o��<`   `   ���<���<���<«�<���<��<���<���<$��<=��<4��<@��<��<@��<4��<=��<$��<���<���<��<���<«�<���<���<`   `   ���<«�<ɫ�<���<���<��<
��<��<M��<���<l��<���<���<���<l��<���<M��<��<
��<��<���<���<ɫ�<«�<`   `   ^��<���<���<���<��<��<���<���<m��<���<���<���<��<���<���<���<m��<���<���<��<��<���<���<���<`   `   ���<���<���<Ы�<*��<��<U��<Ϭ�<n��<���<���<���<��<���<���<���<n��<Ϭ�<U��<��<*��<Ы�<���<���<`   `   ���<���<���<ȫ�<��<���<���<{��<|��<Ĭ�<��<	��<���<	��<��<Ĭ�<|��<{��<���<���<��<ȫ�<���<���<`   `   I��<���<w��<���<	��<��<f��<���<���<ݬ�<��<��<��<��<��<ݬ�<���<���<f��<��<	��<���<w��<���<`   `   ���<���<���<���<
��<��<G��<|��<���<���<���<��<ʬ�<��<���<���<���<|��<G��<��<
��<���<���<���<`   `   ���<���<K��<���<ҫ�<��<!��<>��<���<���<��<��<Ȭ�<��<��<���<���<>��<!��<��<ҫ�<���<K��<���<`   `   `��<M��<0��<X��<~��< ��<���<>��<���<��<���<���<���<���<���<��<���<>��<���< ��<~��<X��<0��<M��<`   `   h��<L��<S��<}��<o��<���<x��<��<]��<Ĭ�<��<��<;��<��<��<Ĭ�<]��<��<x��<���<o��<}��<S��<L��<`   `   t��<8��<G��<���<���<���<8��<3��<3��<g��<w��<���<۬�<���<w��<g��<3��<3��<8��<���<���<���<G��<8��<`   `   _��<��<,��<Q��<c��<���<��<���<N��<K��<���<���<d��<���<���<K��<N��<���<��<���<c��<Q��<,��<��<`   `   ���<Ҫ�<��<1��<[��<���<���<��<	��<C��<���<��<���<��<���<C��<	��<��<���<���<[��<1��<��<Ҫ�<`   `   Ǫ�<���<���<��<\��<���<l��<���<ث�<��<
��<;��<߬�<;��<
��<��<ث�<���<l��<���<\��<��<���<���<`   `   ���<0��<-��<
��<���<x��< ��<��<��<u��<���<��<_��<��<���<u��<��<��< ��<x��<���<
��<-��<0��<`   `   A��<J��<��<��<m��<���<��<���<���<Z��<Q��<r��<O��<r��<Q��<Z��<���<���<��<���<m��<��<��<J��<`   `   ���<G��<���<,��<B��<���<ݭ�<���<���<��<��<7��<\��<7��<��<��<���<���<ݭ�<���<B��<,��<���<G��<`   `   ,��<��<��<\��<[��<���<���<ǭ�<��<���<"��<P��<B��<P��<"��<���<��<ǭ�<���<���<[��<\��<��<��<`   `   "��<^��<{��<y��<���<���<ƭ�<��<��<��<.��<��<˭�<��<.��<��<��<��<ƭ�<���<���<y��<{��<^��<`   `   ���<���<���<���<ȭ�<ƭ�<��<��<��<��<��<��<��<��<��<��<��<��<��<ƭ�<ȭ�<���<���<���<`   `   ��<���<׭�<5��<)��<ʭ�<���<��<��<���<���<��</��<��<���<���<��<��<���<ʭ�<)��<5��<׭�<���<`   `   ��<ڭ�<E��<R��<���<Э�<���<��<��<��<ҭ�<���<ۭ�<���<ҭ�<��<��<��<���<Э�<���<R��<E��<ڭ�<`   `   '��<��<P��<��<���<3��<��<���<��<ޭ�<��<���<���<���<��<ޭ�<��<���<��<3��<���<��<P��<��<`   `   î�<���<���<���<���<���<��<��<P��<��<���<��<ۭ�<��<���<��<P��<��<��<���<���<���<���<���<`   `   !��<��<ޮ�<��<���<���<[��<A��<V��<��<��<��<��<��<��<��<V��<A��<[��<���<���<��<ޮ�<��<`   `   ��<)��<$��<���<Ʈ�<��<���<K��<a��<A��<��<ͭ�<��<ͭ�<��<A��<a��<K��<���<��<Ʈ�<���<$��<)��<`   `   9��<p��<Q��<H��<��<���<t��<M��<O��<V��<)��<��<��<��<)��<V��<O��<M��<t��<���<��<H��<Q��<p��<`   `   ���<���<\��<a��<3��<i��<���<���<.��<���<��<��<ԭ�<��<��<���<.��<���<���<i��<3��<a��<\��<���<`   `   ���<���<���<m��<e��<��<��<���<g��<<��<��<��<���<��<��<<��<g��<���<��<��<e��<m��<���<���<`   `   ��<���<���<���<]��<��<���<���<R��<D��<��<��<׭�<��<��<D��<R��<���<���<��<]��<���<���<���<`   `   _��<���<���<���<Y��<��<ծ�<���<��<��<í�<���<���<���<í�<��<��<���<ծ�<��<Y��<���<���<���<`   `   ��<���<į�<���<a��<��<���<}��<��<3��<��<���<���<���<��<3��<��<}��<���<��<a��<���<į�<���<`   `   ˯�<���<ԯ�<n��<��<��<G��<!��<O��< ��<���<���<^��<���<���< ��<O��<!��<G��<��<��<n��<ԯ�<���<`   `   ���<��<���<;��<���<��<M��<��<��<���<f��<k��<E��<k��<f��<���<��<��<M��<��<���<;��<���<��<`   `   a��<P��<b��<A��<���<���<'��<���<ܭ�<���<���<N��<3��<N��<���<���<ܭ�<���<'��<���<���<A��<b��<P��<`   `   I��<T��<#��<
��<���<&��<��<���<ѭ�<z��<9��<۬�<���<۬�<9��<z��<ѭ�<���<��<&��<���<
��<#��<T��<`   `   ���<��<Ѯ�<ۮ�<���<'��<
��<֭�<���<@��<H��<D��<Y��<D��<H��<@��<���<֭�<
��<'��<���<ۮ�<Ѯ�<��<`   `   C��<��<���<���<r��<G��<(��<���<���<'��<���<���<5��<���<���<'��<���<���<(��<G��<r��<���<���<��<`   `   _��<��<���<u��<��<��< ��<x��<���<
��<-��<0��<���<0��<-��<
��<���<x��< ��<��<��<u��<���<��<`   `   O��<r��<Q��<Z��<���<���<��<���<m��<��<��<J��<A��<J��<��<��<m��<���<��<���<���<Z��<Q��<r��<`   `   \��<7��<��<��<���<���<ݭ�<���<B��<,��<���<G��<���<G��<���<,��<B��<���<ݭ�<���<���<��<��<7��<`   `   B��<P��<"��<���<��<ǭ�<���<���<[��<\��<��<��<,��<��<��<\��<[��<���<���<ǭ�<��<���<"��<P��<`   `   ˭�<��<.��<��<��<��<ƭ�<���<���<y��<{��<^��<"��<^��<{��<y��<���<���<ƭ�<��<��<��<.��<��<`   `   ��<��<��<��<��<��<��<ƭ�<ȭ�<���<���<���<���<���<���<���<ȭ�<ƭ�<��<��<��<��<��<��<`   `   /��<��<���<���<��<��<���<ʭ�<)��<5��<׭�<���<��<���<׭�<5��<)��<ʭ�<���<��<��<���<���<��<`   `   ۭ�<���<ҭ�<��<��<��<���<Э�<���<R��<E��<ڭ�<��<ڭ�<E��<R��<���<Э�<���<��<��<��<ҭ�<���<`   `   ���<���<��<ޭ�<��<���<��<3��<���<��<P��<��<'��<��<P��<��<���<3��<��<���<��<ޭ�<��<���<`   `   ۭ�<��<���<��<P��<��<��<���<���<���<���<���<î�<���<���<���<���<���<��<��<P��<��<���<��<`   `   ��<��<��<��<V��<A��<[��<���<���<��<ޮ�<��<!��<��<ޮ�<��<���<���<[��<A��<V��<��<��<��<`   `   ��<ͭ�<��<A��<a��<K��<���<��<Ʈ�<���<$��<)��<��<)��<$��<���<Ʈ�<��<���<K��<a��<A��<��<ͭ�<`   `   ��<��<)��<V��<O��<M��<t��<���<��<H��<Q��<p��<9��<p��<Q��<H��<��<���<t��<M��<O��<V��<)��<��<`   `   ԭ�<��<��<���<.��<���<���<i��<3��<a��<\��<���<���<���<\��<a��<3��<i��<���<���<.��<���<��<��<`   `   ���<��<��<<��<g��<���<��<��<e��<m��<���<���<���<���<���<m��<e��<��<��<���<g��<<��<��<��<`   `   ׭�<��<��<D��<R��<���<���<��<]��<���<���<���<��<���<���<���<]��<��<���<���<R��<D��<��<��<`   `   ���<���<í�<��<��<���<ծ�<��<Y��<���<���<���<_��<���<���<���<Y��<��<ծ�<���<��<��<í�<���<`   `   ���<���<��<3��<��<}��<���<��<a��<���<į�<���<��<���<į�<���<a��<��<���<}��<��<3��<��<���<`   `   ^��<���<���< ��<O��<!��<G��<��<��<n��<ԯ�<���<˯�<���<ԯ�<n��<��<��<G��<!��<O��< ��<���<���<`   `   E��<k��<f��<���<��<��<M��<��<���<;��<���<��<���<��<���<;��<���<��<M��<��<��<���<f��<k��<`   `   3��<N��<���<���<ܭ�<���<'��<���<���<A��<b��<P��<a��<P��<b��<A��<���<���<'��<���<ܭ�<���<���<N��<`   `   ���<۬�<9��<z��<ѭ�<���<��<&��<���<
��<#��<T��<I��<T��<#��<
��<���<&��<��<���<ѭ�<z��<9��<۬�<`   `   Y��<D��<H��<@��<���<֭�<
��<'��<���<ۮ�<Ѯ�<��<���<��<Ѯ�<ۮ�<���<'��<
��<֭�<���<@��<H��<D��<`   `   5��<���<���<'��<���<���<(��<G��<r��<���<���<��<C��<��<���<���<r��<G��<(��<���<���<'��<���<���<`   `   ���<��<��<j��<ׯ�<���<���<;��<���<��<��<���<��<���<��<��<���<;��<���<���<ׯ�<j��<��<��<`   `   ���<��<W��<k��<���<ʯ�<���<Y��<���<���<���<���<��<���<���<���<���<Y��<���<ʯ�<���<k��<W��<��<`   `   ɮ�<���<n��<|��<���<��<ׯ�<$��<���<���<���<���<��<���<���<���<���<$��<ׯ�<��<���<|��<n��<���<`   `   K��<o��<���<���<���<Я�<¯�<���<R��<z��<���<��<���<��<���<z��<R��<���<¯�<Я�<���<���<���<o��<`   `   ���<̯�<���<���<��<ů�<
��<7��<	��<"��<R��<X��<m��<X��<R��<"��<	��<7��<
��<ů�<��<���<���<̯�<`   `   ���<���<���<���<��<ʯ�<��<��<��<M��<=��<[��<���<[��<=��<M��<��<��<��<ʯ�<��<���<���<���<`   `   J��<���<��<��<��<#��< ��<���<��<���<6��<=��<P��<=��<6��<���<��<���< ��<#��<��<��<��<���<`   `   ���<���<���<Q��<j��<���<���<^��<&��<c��<:��<Q��<-��<Q��<:��<c��<&��<^��<���<���<j��<Q��<���<���<`   `   ��<��<���<���<հ�<���<���<���<M��<J��<9��<J��<)��<J��<9��<J��<M��<���<���<���<հ�<���<���<��<`   `   P��<��<)��<J��<��<���<���<���<n��<k��<j��<G��<F��<G��<j��<k��<n��<���<���<���<��<J��<)��<��<`   `   ��<���<���<t��<��<��<��<˰�<x��<\��<���<>��<T��<>��<���<\��<x��<˰�<��<��<��<t��<���<���<`   `   ��<��<��<|��<l��<���<B��<��<���<[��<F��<��<I��<��<F��<[��<���<��<B��<���<l��<|��<��<��<`   `   ��<S��<5��<��<��<���<��<��<ư�<���<]��<@��<���<@��<]��<���<ư�<��<��<���<��<��<5��<S��<`   `   v��<���<i��<9��<C��<���<���<6��<���<���<d��<,��<��<,��<d��<���<���<6��<���<���<C��<9��<i��<���<`   `   ���<���<���<=��<A��<���<˱�<%��<���<���<O��<"��<د�<"��<O��<���<���<%��<˱�<���<A��<=��<���<���<`   `   ��<���<Ĳ�<J��<��<���<��<���<���<���<?��<?��<W��<?��<?��<���<���<���<��<���<��<J��<Ĳ�<���<`   `   ��<���<Ų�<m��<(��<���<O��<^��<���<��<��<ׯ�<��<ׯ�<��<��<���<^��<O��<���<(��<m��<Ų�<���<`   `   ��<���<���<T��<$��<ر�<z��<9��<o��<=��<��<ݯ�<��<ݯ�<��<=��<o��<9��<z��<ر�<$��<T��<���<���<`   `   ɲ�<���<���<��<ٱ�<���< ��<ܰ�<��<��<ϯ�<��<ǯ�<��<ϯ�<��<��<ܰ�< ��<���<ٱ�<��<���<���<`   `   x��<���<r��<��<߱�<���<��<߰�<e��<ů�<���<���<f��<���<���<ů�<e��<߰�<��<���<߱�<��<r��<���<`   `   P��<B��<3��<���<���<I��<��<���<���<���<Я�<���<n��<���<Я�<���<���<���<��<I��<���<���<3��<B��<`   `   b��<'��<���<���<Z��<���<��<x��<ܯ�<���<���<]��<j��<]��<���<���<ܯ�<x��<��<���<Z��<���<���<'��<`   `   ��<���<E��<h��<C��<��<߰�<��<���<���<H��<��<��<��<H��<���<���<��<߰�<��<C��<h��<E��<���<`   `   L��<˱�<9��<G��<��<���<e��<���<���<}��<��<Ʈ�<Ϯ�<Ʈ�<��<}��<���<���<e��<���<��<G��<9��<˱�<`   `   ��<���<��<��<���<;��<���<���<ׯ�<j��<��<��<���<��<��<j��<ׯ�<���<���<;��<���<��<��<���<`   `   ��<���<���<���<���<Y��<���<ʯ�<���<k��<W��<��<���<��<W��<k��<���<ʯ�<���<Y��<���<���<���<���<`   `   ��<���<���<���<���<$��<ׯ�<��<���<|��<n��<���<ɮ�<���<n��<|��<���<��<ׯ�<$��<���<���<���<���<`   `   ���<��<���<z��<R��<���<¯�<Я�<���<���<���<o��<K��<o��<���<���<���<Я�<¯�<���<R��<z��<���<��<`   `   m��<X��<R��<"��<	��<7��<
��<ů�<��<���<���<̯�<���<̯�<���<���<��<ů�<
��<7��<	��<"��<R��<X��<`   `   ���<[��<=��<M��<��<��<��<ʯ�<��<���<���<���<���<���<���<���<��<ʯ�<��<��<��<M��<=��<[��<`   `   P��<=��<6��<���<��<���< ��<#��<��<��<��<���<J��<���<��<��<��<#��< ��<���<��<���<6��<=��<`   `   -��<Q��<:��<c��<&��<^��<���<���<j��<Q��<���<���<���<���<���<Q��<j��<���<���<^��<&��<c��<:��<Q��<`   `   )��<J��<9��<J��<M��<���<���<���<հ�<���<���<��<��<��<���<���<հ�<���<���<���<M��<J��<9��<J��<`   `   F��<G��<j��<k��<n��<���<���<���<��<J��<)��<��<P��<��<)��<J��<��<���<���<���<n��<k��<j��<G��<`   `   T��<>��<���<\��<x��<˰�<��<��<��<t��<���<���<��<���<���<t��<��<��<��<˰�<x��<\��<���<>��<`   `   I��<��<F��<[��<���<��<B��<���<l��<|��<��<��<��<��<��<|��<l��<���<B��<��<���<[��<F��<��<`   `   ���<@��<]��<���<ư�<��<��<���<��<��<5��<S��<��<S��<5��<��<��<���<��<��<ư�<���<]��<@��<`   `   ��<,��<d��<���<���<6��<���<���<C��<9��<i��<���<v��<���<i��<9��<C��<���<���<6��<���<���<d��<,��<`   `   د�<"��<O��<���<���<%��<˱�<���<A��<=��<���<���<���<���<���<=��<A��<���<˱�<%��<���<���<O��<"��<`   `   W��<?��<?��<���<���<���<��<���<��<J��<Ĳ�<���<��<���<Ĳ�<J��<��<���<��<���<���<���<?��<?��<`   `   ��<ׯ�<��<��<���<^��<O��<���<(��<m��<Ų�<���<��<���<Ų�<m��<(��<���<O��<^��<���<��<��<ׯ�<`   `   ��<ݯ�<��<=��<o��<9��<z��<ر�<$��<T��<���<���<��<���<���<T��<$��<ر�<z��<9��<o��<=��<��<ݯ�<`   `   ǯ�<��<ϯ�<��<��<ܰ�< ��<���<ٱ�<��<���<���<ɲ�<���<���<��<ٱ�<���< ��<ܰ�<��<��<ϯ�<��<`   `   f��<���<���<ů�<e��<߰�<��<���<߱�<��<r��<���<x��<���<r��<��<߱�<���<��<߰�<e��<ů�<���<���<`   `   n��<���<Я�<���<���<���<��<I��<���<���<3��<B��<P��<B��<3��<���<���<I��<��<���<���<���<Я�<���<`   `   j��<]��<���<���<ܯ�<x��<��<���<Z��<���<���<'��<c��<'��<���<���<Z��<���<��<x��<ܯ�<���<���<]��<`   `   ��<��<H��<���<���<��<߰�<��<C��<h��<E��<���<��<���<E��<h��<C��<��<߰�<��<���<���<H��<��<`   `   Ϯ�<Ʈ�<��<}��<���<���<e��<���<��<G��<9��<˱�<L��<˱�<9��<G��<��<���<e��<���<���<}��<��<Ʈ�<`   `   ���<��<N��<S��<���<n��<���<��<c��<���<���<���<��<���<���<���<c��<��<���<n��<���<S��<N��<��<`   `   9��<���<?��<@��<h��<���<��<в�<��<H��<���<}��<���<}��<���<H��<��<в�<��<���<h��<@��<?��<���<`   `   ��<��<P��<m��<���<��<2��<���<���<ڲ�<���<C��<<��<C��<���<ڲ�<���<���<2��<��<���<m��<P��<��<`   `   ���<v��<5��<n��<���<��<X��<q��<y��<���<��<۲�<��<۲�<��<���<y��<q��<X��<��<���<n��<5��<v��<`   `   ���<���<f��<���<��<��<T��<g��<���<���<���<Ҳ�<���<Ҳ�<���<���<���<g��<T��<��<��<���<f��<���<`   `   ��<'��<k��<E��<?��<]��<^��<���<ڲ�<���<ò�<ڲ�<���<ڲ�<ò�<���<ڲ�<���<^��<]��<?��<E��<k��<'��<`   `   Y��<i��<ò�<f��<e��<���<{��<���<Բ�<l��<���<���<��<���<���<l��<Բ�<���<{��<���<e��<f��<ò�<i��<`   `   ���<���<˲�<���<��<²�<v��<���<���<���<���<²�<v��<²�<���<���<���<���<v��<²�<��<���<˲�<���<`   `   \��<���<_��<0��<h��<��<��<ֲ�<���<߲�<y��<���<Ͳ�<���<y��<߲�<���<ֲ�<��<��<h��<0��<_��<���<`   `   ���<��<ݳ�<���<���<���<���<8��<Ҳ�<���<]��<5��<���<5��<]��<���<Ҳ�<8��<���<���<���<���<ݳ�<��<`   `   +��<M��<J��<M��< ��<���<���<;��<���<��<��<���<���<���<��<��<���<;��<���<���< ��<M��<J��<M��<`   `   ��<ȴ�<���<��<c��<ֳ�<��<p��<��<Ҳ�<���<���<���<���<���<Ҳ�<��<p��<��<ֳ�<c��<��<���<ȴ�<`   `   ���<P��<��<��<���<p��<���<���<J��<��<²�<���<���<���<²�<��<J��<���<���<p��<���<��<��<P��<`   `   µ�<y��<u��<��<���<���<���<���<���<M��<в�<���<̲�<���<в�<M��<���<���<���<���<���<��<u��<y��<`   `   ��<���<̵�<���<Ŵ�<���<��<���<���<���<���<���<���<���<���<���<���<���<��<���<Ŵ�<���<̵�<���<`   `   
��<��<��<���<4��<���<R��<ֳ�<i��<���<���<w��<[��<w��<���<���<i��<ֳ�<R��<���<4��<���<��<��<`   `   ���<��<��<n��<3��<��<A��<���<Z��<��<���<[��<C��<[��<���<��<Z��<���<A��<��<3��<n��<��<��<`   `   ڵ�<9��<ֵ�<���<���<[��<��<5��<��<���<H��<*��<-��<*��<H��<���<��<5��<��<[��<���<���<ֵ�<9��<`   `   ��<���<���<���<��<,��<��<I��<Ĳ�<~��<��<��<��<��<��<~��<Ĳ�<I��<��<,��<��<���<���<���<`   `   е�<���<I��<N��<ɴ�<г�<ٳ�<$��<���<���<��<���<���<���<��<���<���<$��<ٳ�<г�<ɴ�<N��<I��<���<`   `   z��<P��<��<���<<��<���<R��<���<\��<F��<s��<C��<q��<C��<s��<F��<\��<���<R��<���<<��<���<��<P��<`   `   ���<���<��<���<��<��<
��<z��<[��<��<T��<T��<W��<T��<T��<��<[��<z��<
��<��<��<���<��<���<`   `   ���<���<д�<A��<���<U��<���<S��<��<���<t��<M��<(��<M��<t��<���<��<S��<���<U��<���<A��<д�<���<`   `   x��<+��<���<ʳ�<O��<ܲ�<���<���<α�<q��<Q��<��<:��<��<Q��<q��<α�<���<���<ܲ�<O��<ʳ�<���<+��<`   `   ��<���<���<���<c��<��<���<n��<���<S��<N��<��<���<��<N��<S��<���<n��<���<��<c��<���<���<���<`   `   ���<|��<���<H��<��<в�<��<���<h��<@��<?��<���<9��<���<?��<@��<h��<���<��<в�<��<H��<���<|��<`   `   <��<C��<���<ڲ�<���<���<2��<��<���<m��<P��<��<��<��<P��<m��<���<��<2��<���<���<ڲ�<���<C��<`   `   ��<۲�<��<���<y��<q��<X��<��<���<n��<5��<v��<���<v��<5��<n��<���<��<X��<q��<y��<���<��<۲�<`   `   ���<Ҳ�<���<���<���<g��<T��<��<��<���<f��<���<���<���<f��<���<��<��<T��<g��<���<���<���<Ҳ�<`   `   ���<ڲ�<ò�<���<ڲ�<���<^��<]��<?��<E��<k��<'��<��<'��<k��<E��<?��<]��<^��<���<ڲ�<���<ò�<ڲ�<`   `   ��<���<���<l��<Բ�<���<{��<���<e��<f��<ò�<i��<Y��<i��<ò�<f��<e��<���<{��<���<Բ�<l��<���<���<`   `   v��<²�<���<���<���<���<v��<²�<��<���<˲�<���<���<���<˲�<���<��<²�<v��<���<���<���<���<²�<`   `   Ͳ�<���<y��<߲�<���<ֲ�<��<��<h��<0��<_��<���<\��<���<_��<0��<h��<��<��<ֲ�<���<߲�<y��<���<`   `   ���<5��<]��<���<Ҳ�<8��<���<���<���<���<ݳ�<��<���<��<ݳ�<���<���<���<���<8��<Ҳ�<���<]��<5��<`   `   ���<���<��<��<���<;��<���<���< ��<M��<J��<M��<+��<M��<J��<M��< ��<���<���<;��<���<��<��<���<`   `   ���<���<���<Ҳ�<��<p��<��<ֳ�<c��<��<���<ȴ�<��<ȴ�<���<��<c��<ֳ�<��<p��<��<Ҳ�<���<���<`   `   ���<���<²�<��<J��<���<���<p��<���<��<��<P��<���<P��<��<��<���<p��<���<���<J��<��<²�<���<`   `   ̲�<���<в�<M��<���<���<���<���<���<��<u��<y��<µ�<y��<u��<��<���<���<���<���<���<M��<в�<���<`   `   ���<���<���<���<���<���<��<���<Ŵ�<���<̵�<���<��<���<̵�<���<Ŵ�<���<��<���<���<���<���<���<`   `   [��<w��<���<���<i��<ֳ�<R��<���<4��<���<��<��<
��<��<��<���<4��<���<R��<ֳ�<i��<���<���<w��<`   `   C��<[��<���<��<Z��<���<A��<��<3��<n��<��<��<���<��<��<n��<3��<��<A��<���<Z��<��<���<[��<`   `   -��<*��<H��<���<��<5��<��<[��<���<���<ֵ�<9��<ڵ�<9��<ֵ�<���<���<[��<��<5��<��<���<H��<*��<`   `   ��<��<��<~��<Ĳ�<I��<��<,��<��<���<���<���<��<���<���<���<��<,��<��<I��<Ĳ�<~��<��<��<`   `   ���<���<��<���<���<$��<ٳ�<г�<ɴ�<N��<I��<���<е�<���<I��<N��<ɴ�<г�<ٳ�<$��<���<���<��<���<`   `   q��<C��<s��<F��<\��<���<R��<���<<��<���<��<P��<z��<P��<��<���<<��<���<R��<���<\��<F��<s��<C��<`   `   W��<T��<T��<��<[��<z��<
��<��<��<���<��<���<���<���<��<���<��<��<
��<z��<[��<��<T��<T��<`   `   (��<M��<t��<���<��<S��<���<U��<���<A��<д�<���<���<���<д�<A��<���<U��<���<S��<��<���<t��<M��<`   `   :��<��<Q��<q��<α�<���<���<ܲ�<O��<ʳ�<���<+��<x��<+��<���<ʳ�<O��<ܲ�<���<���<α�<q��<Q��<��<`   `   c��<���<��<���<���<&��<ô�<p��<���<3��<���<���<���<���<���<3��<���<p��<ô�<&��<���<���<��<���<`   `   ���<���<в�<P��<г�<��<n��<ݴ�<%��<���<��<)��<~��<)��<��<���<%��<ݴ�<n��<��<г�<P��<в�<���<`   `   ��</��<��<x��<��<��<p��<��<E��<Q��<l��<���<��<���<l��<Q��<E��<��<p��<��<��<x��<��</��<`   `   ��<h��<���<��<���<ܳ�<\��<���<M��<J��<E��<���<͵�<���<E��<J��<M��<���<\��<ܳ�<���<��<���<h��<`   `   c��<���<���<��<���<1��<^��<W��<��<$��<"��<.��<E��<.��<"��<$��<��<W��<^��<1��<���<��<���<���<`   `   ^��<-��< ��<A��<\��<{��<v��<v��<���<Ӵ�<��<��<��<��<��<Ӵ�<���<v��<v��<{��<\��<A��< ��<-��<`   `   ��<���<���<˴�<���<ش�<��<ܴ�<���<���<��<��<0��<��<��<���<���<ܴ�<��<ش�<���<˴�<���<���<`   `   ���<J��<M��<���<F��<6��<X��<*��<��<��<��<��<ݴ�<��<��<��<��<*��<X��<6��<F��<���<M��<J��<`   `   ��<��<��<��<���<^��<l��<=��<6��<��<,��<��<ô�<��<,��<��<6��<=��<l��<^��<���<��<��<��<`   `   ���<��<���<R��<:��<��<׵�<l��<U��<��<
��<)��<��<)��<
��<��<U��<l��<׵�<��<:��<R��<���<��<`   `   ���<���<E��<��<���<���<%��<���<ε�<!��<ܴ�<��<��<��<ܴ�<!��<ε�<���<%��<���<���<��<E��<���<`   `   ��<
��<з�<���<Q��<ն�<���<!��<���<}��<��<��<̴�<��<��<}��<���<!��<���<ն�<Q��<���<з�<
��<`   `   ���<���<x��<��<���<W��<��<d��<���<c��<2��<��<���<��<2��<c��<���<d��<��<W��<���<��<x��<���<`   `   ��<��<���<���<:��<·�<��<j��<ŵ�<W��<%��<��<д�<��<%��<W��<ŵ�<j��<��<·�<:��<���<���<��<`   `   ���<E��<���<���<g��<���<��<���<���<a��<>��<��<���<��<>��<a��<���<���<��<���<g��<���<���<E��<`   `   ݹ�<���<���<���<Z��<���<Y��<���<���<4��<9��<���<k��<���<9��<4��<���<���<Y��<���<Z��<���<���<���<`   `   ���<ȹ�<��<��<`��<���<��</��<���<��<��<~��<n��<~��<��<��<���</��<��<���<`��<��<��<ȹ�<`   `   ���<̹�<��<޸�<'��<���<���<)��<��<��<���<K��<%��<K��<���<��<��<)��<���<���<'��<޸�<��<̹�<`   `   (��<I��<Ը�<���<���<���<��<	��<���<���<f��<���<���<���<f��<���<���<	��<��<���<���<���<Ը�<I��<`   `   ڸ�< ��<ĸ�<J��<ҷ�<0��<b��<���<��<h��<��<��<��<��<��<h��<��<���<b��<0��<ҷ�<J��<ĸ�< ��<`   `   ��<ʸ�<t��<۷�<��<׶�<��<t��<���<��<���<���<���<���<���<��<���<t��<��<׶�<��<۷�<t��<ʸ�<`   `   ���<��<��<n��<��<���<���<L��<���<���<��<V��<���<V��<��<���<���<L��<���<���<��<n��<��<��<`   `   ��<���<���<��<���<��<��<ʴ�<��<d��<F��<*��<���<*��<F��<d��<��<ʴ�<��<��<���<��<���<���<`   `   p��<��<��<x��<1��<��<���<w��<���<k��<��<���<���<���<��<k��<���<w��<���<��<1��<x��<��<��<`   `   ���<���<���<3��<���<p��<´�<&��<���<���<��<���<c��<���<��<���<���<&��<´�<p��<���<3��<���<���<`   `   ~��<)��<��<���<%��<ݴ�<n��<��<г�<P��<в�<���<���<���<в�<P��<г�<��<n��<ݴ�<%��<���<��<)��<`   `   ��<���<l��<Q��<E��<��<p��<��<��<x��<��</��<��</��<��<x��<��<��<p��<��<E��<Q��<l��<���<`   `   ͵�<���<E��<J��<M��<���<\��<ܳ�<���<��<���<h��<��<h��<���<��<���<ܳ�<\��<���<M��<J��<E��<���<`   `   E��<.��<"��<$��<��<W��<^��<1��<���<��<���<���<c��<���<���<��<���<1��<^��<W��<��<$��<"��<.��<`   `   ��<��<��<Ӵ�<���<v��<v��<{��<\��<A��< ��<-��<^��<-��< ��<A��<\��<{��<v��<v��<���<Ӵ�<��<��<`   `   0��<��<��<���<���<ܴ�<��<ش�<���<˴�<���<���<��<���<���<˴�<���<ش�<��<ܴ�<���<���<��<��<`   `   ݴ�<��<��<��<��<*��<X��<6��<F��<���<M��<J��<���<J��<M��<���<F��<6��<X��<*��<��<��<��<��<`   `   ô�<��<,��<��<6��<=��<l��<^��<���<��<��<��<��<��<��<��<���<^��<l��<=��<6��<��<,��<��<`   `   ��<)��<
��<��<U��<l��<׵�<��<:��<R��<���<��<���<��<���<R��<:��<��<׵�<l��<U��<��<
��<)��<`   `   ��<��<ܴ�<!��<ε�<���<%��<���<���<��<E��<���<���<���<E��<��<���<���<%��<���<ε�<!��<ܴ�<��<`   `   ̴�<��<��<}��<���<!��<���<ն�<Q��<���<з�<
��<��<
��<з�<���<Q��<ն�<���<!��<���<}��<��<��<`   `   ���<��<2��<c��<���<d��<��<W��<���<��<x��<���<���<���<x��<��<���<W��<��<d��<���<c��<2��<��<`   `   д�<��<%��<W��<ŵ�<j��<��<·�<:��<���<���<��<��<��<���<���<:��<·�<��<j��<ŵ�<W��<%��<��<`   `   ���<��<>��<a��<���<���<��<���<g��<���<���<E��<���<E��<���<���<g��<���<��<���<���<a��<>��<��<`   `   k��<���<9��<4��<���<���<Y��<���<Z��<���<���<���<ݹ�<���<���<���<Z��<���<Y��<���<���<4��<9��<���<`   `   n��<~��<��<��<���</��<��<���<`��<��<��<ȹ�<���<ȹ�<��<��<`��<���<��</��<���<��<��<~��<`   `   %��<K��<���<��<��<)��<���<���<'��<޸�<��<̹�<���<̹�<��<޸�<'��<���<���<)��<��<��<���<K��<`   `   ���<���<f��<���<���<	��<��<���<���<���<Ը�<I��<(��<I��<Ը�<���<���<���<��<	��<���<���<f��<���<`   `   ��<��<��<h��<��<���<b��<0��<ҷ�<J��<ĸ�< ��<ڸ�< ��<ĸ�<J��<ҷ�<0��<b��<���<��<h��<��<��<`   `   ���<���<���<��<���<t��<��<׶�<��<۷�<t��<ʸ�<��<ʸ�<t��<۷�<��<׶�<��<t��<���<��<���<���<`   `   ���<V��<��<���<���<L��<���<���<��<n��<��<��<���<��<��<n��<��<���<���<L��<���<���<��<V��<`   `   ���<*��<F��<d��<��<ʴ�<��<��<���<��<���<���<��<���<���<��<���<��<��<ʴ�<��<d��<F��<*��<`   `   ���<���<��<k��<���<w��<���<��<1��<x��<��<��<p��<��<��<x��<1��<��<���<w��<���<k��<��<���<`   `   J��<���<���<��<���<��<޶�<p��<M��<Ѹ�<`��<���<���<���<`��<Ѹ�<M��<p��<޶�<��<���<��<���<���<`   `   Y��<ٴ�<���<��<���<��<���<<��<��<���<���<��<��<��<���<���<��<<��<���<��<���<��<���<ٴ�<`   `   Z��<���<���<��<���<���<���<��<ȷ�<,��<9��<���<@��<���<9��<,��<ȷ�<��<���<���<���<��<���<���<`   `   ���<��<)��<K��<���<*��<���<���<"��<���<��<G��<��<G��<��<���<"��<���<���<*��<���<K��<)��<��<`   `   µ�<ӵ�<ҵ�<���<��<���<��<8��<��<2��<���<���<���<���<���<2��<��<8��<��<���<��<���<ҵ�<ӵ�<`   `   ��<:��<+��<H��<���<���<��<^��<4��<h��<f��<.��<��<.��<f��<h��<4��<^��<��<���<���<H��<+��<:��<`   `   z��<��<��<���<	��<��<���<
��<9��<���<u��<6��<���<6��<u��<���<9��<
��<���<��<	��<���<��<��<`   `   ��<'��<ڷ�<���<���<ҷ�<���<H��<Z��<p��<��<ڶ�<K��<ڶ�<��<p��<Z��<H��<���<ҷ�<���<���<ڷ�<'��<`   `   ɸ�<���<���<���<T��<u��<��<ٷ�<���<<��<B��<��<��<��<B��<<��<���<ٷ�<��<u��<T��<���<���<���<`   `   ���<`��<}��<���<��<���<D��<I��<��<~��<���<g��<��<g��<���<~��<��<I��<D��<���<��<���<}��<`��<`   `   ���<���<|��<)��<���<\��<���<���<��<���<u��<7��<���<7��<u��<���<��<���<���<\��<���<)��<|��<���<`   `   @��<f��<9��<���<n��<���<���<���<&��< ��<l��<c��<t��<c��<l��< ��<&��<���<���<���<n��<���<9��<f��<`   `   ��<D��<���<V��<��<��<���<��<z��<I��<���<���<���<���<���<I��<z��<��<���<��<��<V��<���<D��<`   `   ��<���<|��<���<���<���<׹�<k��<���<��<}��<8��<+��<8��<}��<��<���<k��<׹�<���<���<���<|��<���<`   `   "��<X��<��<��<ƻ�<$��<:��<k��<���<'��<|��<��<:��<��<|��<'��<���<k��<:��<$��<ƻ�<��<��<X��<`   `   =��<���<U��<���<ʻ�<���<��<6��<���<8��<Q��<��<L��<��<Q��<8��<���<6��<��<���<ʻ�<���<U��<���<`   `   P��<}��<H��<��<���<���<��<>��<w��<���<��<���<��<���<��<���<w��<>��<��<���<���<��<H��<}��<`   `   ���<]��<��<ü�<���<
��<���<��<��<'��<��<r��<���<r��<��<'��<��<��<���<
��<���<ü�<��<]��<`   `   ���<M��<���<,��</��<���<E��<���<���<���<���<���<��<���<���<���<���<���<E��<���</��<,��<���<M��<`   `   ��<ټ�<���<���<���<K��<��<a��<���<u��<���<z��<z��<z��<���<u��<���<a��<��<K��<���<���<���<ټ�<`   `   ��<��<���<e��<���<���<ø�<���<���<H��<���<S��<��<S��<���<H��<���<���<ø�<���<���<e��<���<��<`   `   ɻ�<}��<��<Ϻ�<��<���<e��<>��<6��<��<o��<��<���<��<o��<��<6��<>��<e��<���<��<Ϻ�<��<}��<`   `   1��<���<���<&��<���<p��<	��<��<%��<Ƶ�<���<���<���<���<���<Ƶ�<%��<��<	��<p��<���<&��<���<���<`   `   ��<:��<��<k��<	��<��<W��<���<
��<l��<^��<���<���<���<^��<l��<
��<���<W��<��<	��<k��<��<:��<`   `   ���<���<`��<Ѹ�<M��<p��<޶�<��<���<��<���<���<J��<���<���<��<���<��<޶�<p��<M��<Ѹ�<`��<���<`   `   ��<��<���<���<��<<��<���<��<���<��<���<ٴ�<Y��<ٴ�<���<��<���<��<���<<��<��<���<���<��<`   `   @��<���<9��<,��<ȷ�<��<���<���<���<��<���<���<Z��<���<���<��<���<���<���<��<ȷ�<,��<9��<���<`   `   ��<G��<��<���<"��<���<���<*��<���<K��<(��<��<���<��<(��<K��<���<*��<���<���<"��<���<��<G��<`   `   ���<���<���<2��<��<8��<��<���<��<���<ҵ�<ӵ�<µ�<ӵ�<ҵ�<���<��<���<��<8��<��<2��<���<���<`   `   ��<.��<f��<h��<4��<^��<��<���<���<H��<+��<:��<��<:��<+��<H��<���<���<��<^��<4��<h��<f��<.��<`   `   ���<6��<u��<���<9��<
��<���<��<	��<���<��<��<z��<��<��<���<	��<��<���<
��<9��<���<u��<6��<`   `   K��<ڶ�<��<p��<Z��<H��<���<ҷ�<���<���<ڷ�<'��<��<'��<ڷ�<���<���<ҷ�<���<H��<Z��<p��<��<ڶ�<`   `   ��<��<B��<<��<���<ٷ�<��<u��<T��<���<���<���<ɸ�<���<���<���<T��<u��<��<ٷ�<���<<��<B��<��<`   `   ��<g��<���<~��<��<I��<D��<���<��<���<}��<`��<���<`��<}��<���<��<���<D��<I��<��<~��<���<g��<`   `   ���<7��<u��<���<��<���<���<\��<���<)��<|��<���<���<���<|��<)��<���<\��<���<���<��<���<u��<7��<`   `   t��<c��<l��< ��<&��<���<���<���<n��<���<9��<f��<@��<f��<9��<���<n��<���<���<���<&��< ��<l��<c��<`   `   ���<���<���<I��<z��<��<���<��<��<V��<���<D��<��<D��<���<V��<��<��<���<��<z��<I��<���<���<`   `   +��<8��<}��<��<���<k��<׹�<���<���<���<|��<���<��<���<|��<���<���<���<׹�<k��<���<��<}��<8��<`   `   :��<��<|��<'��<���<k��<:��<$��<ƻ�<��<��<X��<"��<X��<��<��<ƻ�<$��<:��<k��<���<'��<|��<��<`   `   L��<��<Q��<8��<���<6��<��<���<ʻ�<���<U��<���<=��<���<U��<���<ʻ�<���<��<6��<���<8��<Q��<��<`   `   ��<���<��<���<w��<>��<��<���<���<��<H��<}��<P��<}��<H��<��<���<���<��<>��<w��<���<��<���<`   `   ���<r��<��<'��<��<��<���<
��<���<ü�<��<]��<���<]��<��<ü�<���<
��<���<��<��<'��<��<r��<`   `   ��<���<���<���<���<���<E��<���</��<,��<���<M��<���<M��<���<,��</��<���<E��<���<���<���<���<���<`   `   z��<z��<���<u��<���<a��<��<K��<���<���<���<ټ�<��<ټ�<���<���<���<K��<��<a��<���<u��<���<z��<`   `   ��<S��<���<H��<���<���<ø�<���<���<e��<���<��<��<��<���<e��<���<���<ø�<���<���<H��<���<S��<`   `   ���<��<o��<��<6��<>��<e��<���<��<Ϻ�<��<}��<ɻ�<}��<��<Ϻ�<��<���<e��<>��<6��<��<o��<��<`   `   ���<���<���<Ƶ�<%��<��<	��<p��<���<&��<���<���<1��<���<���<&��<���<p��<	��<��<%��<Ƶ�<���<���<`   `   ���<���<^��<l��<
��<���<W��<��<	��<k��<��<:��<��<:��<��<k��<	��<��<W��<���<
��<l��<^��<���<`   `   #��<���<��<8��<C��<c��<Q��<(��<��<���<5��<¼�<ռ�<¼�<5��<���<��<(��<Q��<c��<C��<8��<��<���<`   `   p��<���<��<���<'��<ݷ�<���<���<j��<���<|��<
��<���<
��<|��<���<j��<���<���<ݷ�<'��<���<��<���<`   `   /��<��<t��<���<8��<���<���<D��<���<V��<��<G��<&��<G��<��<V��<���<D��<���<���<8��<���<t��<��<`   `   ¶�<K��<���<��<���<��<Z��<.��<x��<���<H��<k��<n��<k��<H��<���<x��<.��<Z��<��<���<��<���<K��<`   `   F��< ��<U��<q��<з�<��<,��<��<{��<ڹ�<���</��<r��</��<���<ڹ�<{��<��<,��<��<з�<q��<U��< ��<`   `    ��<��<K��<c��<}��<���<ĸ�<��<J��<a��<���<չ�<��<չ�<���<a��<J��<��<ĸ�<���<}��<c��<K��<��<`   `   ���<M��<I��<t��<���<i��<q��<y��<n��<(��<}��<���<2��<���<}��<(��<n��<y��<q��<i��<���<t��<I��<M��<`   `    ��<k��<>��<��<��<Ϲ�<���<ι�<���<g��<���<���<���<���<���<g��<���<ι�<���<Ϲ�<��<��<>��<k��<`   `   ���<���<q��<'��<��<Ժ�<L��<1��<��<���<���<���<���<���<���<���<��<1��<L��<Ժ�<��<'��<q��<���<`   `   9��<ݼ�<���<w��<��<���<��<Ⱥ�<5��< ��<���<6��<¹�<6��<���< ��<5��<Ⱥ�<��<���<��<w��<���<ݼ�<`   `   V��<���<ѽ�<i��<Ӽ�<K��<һ�<T��<x��<_��<��<���<���<���<��<_��<x��<T��<һ�<K��<Ӽ�<i��<ѽ�<���<`   `   [��<%��<���<���<��<<��<v��<���<ú�<L��<ع�<���<{��<���<ع�<L��<ú�<���<v��<<��<��<���<���<%��<`   `   t��<��<Կ�<���<׾�<н�<��<��<W��<z��<ѹ�<���<6��<���<ѹ�<z��<W��<��<��<н�<׾�<���<Կ�<��<`   `   @��<���<���<��<��<1��<_��<X��<l��<��<���<���<H��<���<���<��<l��<X��<_��<1��<��<��<���<���<`   `   ���<S��<<��<���<���<���<���<>��<<��<M��<ù�<���<,��<���<ù�<M��<<��<>��<���<���<���<���<<��<S��<`   `   <��<���<���<���<���<��<���<R��<R��<0��<���<B��<Ҹ�<B��<���<0��<R��<R��<���<��<���<���<���<���<`   `   ���<)��<i��<b��<ǿ�<ž�<x��<V��<��<��<`��<͸�<E��<͸�<`��<��<��<V��<x��<ž�<ǿ�<b��<i��<)��<`   `   !��<���<[��<u��<���<^��<"��<��<o��<��<��<5��<��<5��<��<��<o��<��<"��<^��<���<u��<[��<���<`   `   ���<K��<��<���<[��<��<���<���<��<���<x��<ŷ�<��<ŷ�<x��<���<��<���<���<��<[��<���<��<K��<`   `   q��<���<6��<���<���<���<V��<��<���<ڸ�<ݷ�<C��<b��<C��<ݷ�<ڸ�<���<��<V��<���<���<���<6��<���<`   `   z��<`��<���<��< ��<��<���<#��<3��<��<B��<׶�<���<׶�<B��<��<3��<#��<���<��< ��<��<���<`��<`   `   a��<���<'��<;��<K��<3��<��<d��<���<���<���<P��<`��<P��<���<���<���<d��<��<3��<K��<;��<'��<���<`   `   ���<���<+��<g��<���<t��<w��<��<��<@��<n��<��<ǵ�<��<n��<@��<��<��<w��<t��<���<g��<+��<���<`   `   ҽ�<���<3��<���<���<���<���<���<���<���<_��<ѵ�<^��<ѵ�<_��<���<���<���<���<���<���<���<3��<���<`   `   ռ�<¼�<4��<���<��<(��<Q��<c��<C��<8��<��<���<#��<���<��<8��<C��<c��<Q��<(��<��<���<4��<¼�<`   `   ���<
��<|��<���<j��<���<���<ݷ�<'��<���<��<���<p��<���<��<���<'��<ݷ�<���<���<j��<���<|��<
��<`   `   &��<F��<��<V��<���<D��<���<���<8��<���<t��<��</��<��<t��<���<8��<���<���<D��<���<V��<��<F��<`   `   n��<k��<H��<���<x��<.��<Z��<��<���<��<���<K��<¶�<K��<���<��<���<��<Z��<.��<x��<���<H��<k��<`   `   r��</��<���<ڹ�<{��<��<,��<��<з�<q��<U��< ��<F��< ��<U��<q��<з�<��<,��<��<{��<ڹ�<���</��<`   `   ��<չ�<���<a��<J��<��<ĸ�<���<}��<c��<K��<��< ��<��<K��<c��<}��<���<ĸ�<��<J��<a��<���<չ�<`   `   2��<���<}��<(��<n��<y��<q��<i��<���<t��<I��<M��<���<M��<I��<t��<���<i��<q��<y��<n��<(��<}��<���<`   `   ���<���<���<g��<���<ι�<���<Ϲ�<��<��<>��<k��< ��<k��<>��<��<��<Ϲ�<���<ι�<���<g��<���<���<`   `   ���<���<���<���<��<1��<L��<Ժ�<��<'��<q��<���<���<���<q��<'��<��<Ժ�<L��<1��<��<���<���<���<`   `   ¹�<6��<���< ��<5��<Ⱥ�<��<���<��<w��<���<ݼ�<9��<ݼ�<���<w��<��<���<��<Ⱥ�<5��< ��<���<6��<`   `   ���<���<��<_��<x��<T��<һ�<K��<Ӽ�<i��<ѽ�<���<V��<���<ѽ�<i��<Ӽ�<K��<һ�<T��<x��<_��<��<���<`   `   {��<���<ع�<L��<ú�<���<v��<<��<��<���<���<%��<[��<%��<���<���<��<<��<v��<���<ú�<L��<ع�<���<`   `   6��<���<ѹ�<z��<W��<��<��<н�<׾�<���<Կ�<��<t��<��<Կ�<���<׾�<н�<��<��<W��<z��<ѹ�<���<`   `   H��<���<���<��<l��<X��<_��<1��<��<��<���<���<@��<���<���<��<��<1��<_��<X��<l��<��<���<���<`   `   ,��<���<ù�<M��<<��<>��<���<���<���<���<<��<S��<���<S��<<��<���<���<���<���<>��<<��<M��<ù�<���<`   `   Ҹ�<B��<���<0��<R��<R��<���<��<���<���<���<���<<��<���<���<���<���<��<���<R��<R��<0��<���<B��<`   `   E��<͸�<`��<��<��<V��<x��<ž�<ǿ�<b��<i��<)��<���<)��<i��<b��<ǿ�<ž�<x��<V��<��<��<`��<͸�<`   `   ��<5��<��<��<o��<��<"��<^��<���<u��<[��<���<!��<���<[��<u��<���<^��<"��<��<o��<��<��<5��<`   `   ��<ŷ�<x��<���<��<���<���<��<[��<���<��<K��<���<K��<��<���<[��<��<���<���<��<���<x��<ŷ�<`   `   b��<C��<ݷ�<ڸ�<���<��<W��<���<���<���<6��<���<q��<���<6��<���<���<���<W��<��<���<ڸ�<ݷ�<C��<`   `   ���<׶�<B��<��<3��<#��<���<��< ��<��<���<`��<z��<`��<���<��< ��<��<���<#��<3��<��<B��<׶�<`   `   a��<P��<���<���<���<d��<��<3��<K��<;��<'��<���<a��<���<'��<;��<K��<3��<��<d��<���<���<���<P��<`   `   ǵ�<��<o��<@��<��<��<w��<t��<���<g��<+��<���<���<���<+��<g��<���<t��<w��<��<��<@��<o��<��<`   `   ^��<ѵ�<_��<���<���<���<���<���<���<���<3��<���<ҽ�<���<3��<���<���<���<���<���<���<���<_��<ѵ�<`   `   ƶ�<j��<��<��<���<��<��<���<���<��<���<߿�<?��<߿�<���<��<���<���<��<��<���<��<��<j��<`   `   ���<P��<��<η�<���<���<[��<���<ͼ�<ֽ�<���<���<پ�<���<���<ֽ�<ͼ�<���<[��<���<���<η�<��<P��<`   `   ���<ض�<g��<���<w��<���<O��<c��<4��<"��<���<��<k��<��<���<"��<4��<c��<O��<���<w��<���<g��<ض�<`   `   ���<���<��<9��<��<޹�<���<���<��<���<���<��<k��<��<���<���<��<���<���<޹�<��<9��<��<���<`   `   a��<_��<��<B��<���<���<���<���<t��<-��<;��<b��<��<b��<;��<-��<t��<���<���<���<���<B��<��<_��<`   `   ��<���<ι�<���<���<̺�<0��<Ӻ�<r��<޻�<���<<��<���<<��<���<޻�<r��<Ӻ�<0��<̺�<���<���<ι�<���<`   `   λ�<K��<Ժ�<��<��<x��<ֻ�<|��<һ�<���<���<��<h��<��<���<���<һ�<|��<ֻ�<x��<��<��<Ժ�<K��<`   `   ���<���<���<Լ�<���<��<C��<%��<��<ֻ�<ݻ�<���<3��<���<ݻ�<ֻ�<��<%��<C��<��<���<Լ�<���<���<`   `   m��<y��<p��<,��<ʽ�<n��<>��<���<J��<6��<��<}��<@��<}��<��<6��<J��<���<>��<n��<ʽ�<,��<p��<y��<`   `   4��<*��<��<R��<
��<���<��<:��<���<L��<���<���<���<���<���<L��<���<:��<��<���<
��<R��<��<*��<`   `   ���<���<i��<���<z��<���<���<��<Q��<���<��<���<һ�<���<��<���<Q��<��<���<���<z��<���<i��<���<`   `   ���<i��<���<#��<V��<w��<]��<���<��<Ҽ�<\��<��<���<��<\��<Ҽ�<��<���<]��<w��<V��<#��<���<i��<`   `   ���<���<*��<C��<.��<���<G��<��<��<��<S��<��<���<��<S��<��<��<��<G��<���<.��<C��<*��<���<`   `   ��<���<O��<���<1��<H��<���<A��<��<-��<u��<��<ֻ�<��<u��<-��<��<A��<���<H��<1��<���<O��<���<`   `   &��<���<���<'��<���<I��<���<���<W��<:��<5��<x��<9��<x��<5��<:��<W��<���<���<I��<���<'��<���<���<`   `   Q��<���<A��<���<1��<w��<��<���<8��<ʼ�<ػ�<e��<̺�<e��<ػ�<ʼ�<8��<���<��<w��<1��<���<A��<���<`   `   j��<��<���<���<J��<~��<���<6��<���<L��<p��<K��<���<K��<p��<L��<���<6��<���<~��<J��<���<���<��<`   `   ��<��<���<$��<��<:��<���<Ѿ�<]��<��<l��<R��<۹�<R��<l��<��<]��<Ѿ�<���<:��<��<$��<���<��<`   `   ���<���<��<���<y��<���<*��<Z��<���<4��<���<���<l��<���<���<4��<���<Z��<*��<���<y��<���<��<���<`   `   ���<���<��<��<��<���<a��<W��<���<M��<���<���<a��<���<���<M��<���<W��<a��<���<��<��<��<���<`   `   ���<���<'��<9��<���<��<i��<���<7��<���<��<?��<���<?��<��<���<7��<���<i��<��<���<9��<'��<���<`   `   ���<���<���<���<���<c��<x��<C��<��<��<5��<���<{��<���<5��<��<��<C��<x��<c��<���<���<���<���<`   `   ���<9��<���<���<���<\��<q��<=��<ù�<;��<ķ�<ն�<���<ն�<ķ�<;��<ù�<=��<q��<\��<���<���<���<9��<`   `   ���<&��<���<���<v��<h��<���<S��<��<���<���<���<b��<���<���<���<��<S��<���<h��<v��<���<���<&��<`   `   ?��<߿�<���<��<���<���<��<��<���<��<��<j��<ƶ�<j��<��<��<���<��<��<���<���<��<���<߿�<`   `   پ�<���<���<ֽ�<ͼ�<���<[��<���<���<η�<��<P��<���<P��<��<η�<���<���<[��<���<ͼ�<ֽ�<���<���<`   `   k��<��<���<"��<4��<c��<O��<���<w��<���<g��<ض�<���<ض�<g��<���<w��<���<O��<c��<4��<"��<���<��<`   `   k��<��<���<���<��<���<���<޹�<��<9��<��<���<���<���<��<9��<��<޹�<���<���<��<���<���<��<`   `   ��<b��<;��<-��<t��<���<���<���<���<B��<��<_��<a��<_��<��<B��<���<���<���<���<t��<-��<;��<b��<`   `   ���<<��<���<޻�<r��<Ӻ�<0��<̺�<���<���<ι�<���<��<���<ι�<���<���<̺�<0��<Ӻ�<r��<޻�<���<<��<`   `   g��<��<���<���<һ�<|��<ֻ�<x��<��<��<Ժ�<K��<λ�<K��<Ժ�<��<��<x��<ֻ�<|��<һ�<���<���<��<`   `   3��<���<ݻ�<ֻ�<��<%��<C��<��<���<Լ�<���<���<���<���<���<Լ�<���<��<C��<%��<��<ֻ�<ݻ�<���<`   `   @��<}��<��<6��<J��<���<>��<n��<ʽ�<,��<p��<y��<m��<y��<p��<,��<ʽ�<n��<>��<���<J��<6��<��<}��<`   `   ���<���<���<L��<���<:��<��<���<
��<R��<��<*��<4��<*��<��<R��<
��<���<��<:��<���<L��<���<���<`   `   һ�<���<��<���<Q��<��<���<���<z��<���<i��<���<���<���<i��<���<z��<���<���<��<Q��<���<��<���<`   `   ���<��<\��<Ҽ�<��<���<]��<w��<V��<#��<���<i��<���<i��<���<#��<V��<w��<]��<���<��<Ҽ�<\��<��<`   `   ���<��<S��<��<��<��<G��<���<.��<C��<*��<���<���<���<*��<C��<.��<���<G��<��<��<��<S��<��<`   `   ֻ�<��<u��<-��<��<A��<���<H��<1��<���<O��<���<��<���<O��<���<1��<H��<���<A��<��<-��<u��<��<`   `   9��<x��<5��<:��<W��<���<���<I��<���<'��<���<���<&��<���<���<'��<���<I��<���<���<W��<:��<5��<x��<`   `   ̺�<e��<ػ�<ʼ�<8��<���<��<w��<1��<���<A��<���<Q��<���<A��<���<1��<w��<��<���<8��<ʼ�<ػ�<e��<`   `   ���<K��<p��<L��<���<6��<���<~��<J��<���<���<��<j��<��<���<���<J��<~��<���<6��<���<L��<p��<K��<`   `   ۹�<R��<l��<��<]��<Ѿ�<���<:��<��<$��<���<��<��<��<���<$��<��<:��<���<Ѿ�<]��<��<l��<R��<`   `   l��<���<���<4��<���<Z��<*��<���<y��<���<��<���<���<���<��<���<y��<���<*��<Z��<���<4��<���<���<`   `   a��<���<���<M��<���<W��<a��<���<��<��<��<���<���<���<��<��<��<���<a��<W��<���<M��<���<���<`   `   ���<?��<��<���<7��<���<i��<��<���<9��<'��<���<���<���<'��<9��<���<��<i��<���<7��<���<��<?��<`   `   {��<���<5��<��<��<C��<x��<c��<���<���<���<���<���<���<���<���<���<c��<x��<C��<��<��<5��<���<`   `   ���<ն�<ķ�<;��<ù�<=��<q��<\��<���<���<���<9��<���<9��<���<���<���<\��<q��<=��<ù�<;��<ķ�<ն�<`   `   b��<���<���<���<��<S��<���<h��<v��<���<���<&��<���<&��<���<���<v��<h��<���<S��<��<���<���<���<`   `   ���<���<4��<e��<���<P��<C��<��<U��<���<���<���<���<���<���<���<U��<��<C��<P��<���<e��<4��<���<`   `   ���<��<���<>��<I��<��<���<
��<���<a��<o��<��</��<��<o��<a��<���<
��<���<��<I��<>��<���<��<`   `   ���<[��<��<{��<���<���<��<��<���<���<C��<���<���<���<C��<���<���<��<��<���<���<{��<��<[��<`   `   ��<V��<q��<��<��<���<���<���<���<���<e��<ο�<¿�<ο�<e��<���<���<���<���<���<��<��<q��<V��<`   `   ���<���<���<=��<���<3��<7��<���<@��<���<���<��<���<��<���<���<@��<���<7��<3��<���<=��<���<���<`   `   ɺ�<��<u��<���<)��<6��<���<\��<���<ν�<���</��<��</��<���<ν�<���<\��<���<6��<)��<���<u��<��<`   `   ���<��<i��<B��<F��< ��<��<T��<���<���<���<��<s��<��<���<���<���<T��<��< ��<F��<B��<i��<��<`   `   '��<-��<I��<��<���<¾�<Z��<��<���<ý�<^��<���<��<���<^��<ý�<���<��<Z��<¾�<���<��<I��<-��<`   `   ���<k��</��<���<x��<��<���<��<���<��<̽�<ܽ�<���<ܽ�<̽�<��<���<��<���<��<x��<���</��<k��<`   `   ���<���<f��<���<&��<5��<���<ݿ�<b��<���<4��<<��<���<<��<4��<���<b��<ݿ�<���<5��<&��<���<f��<���<`   `   ��<��<���<&��<O��<
��<��<���<̿�<̾�<'��<׽�<L��<׽�<'��<̾�<̿�<���<��<
��<O��<&��<���<��<`   `   f��<@��<���<���<���<]��<+��<���<N��<Z��<{��<ݽ�<���<ݽ�<{��<Z��<N��<���<+��<]��<���<���<���<@��<`   `   ���<���<(��<e��<��<q��<���<H��<���<���<���<ٽ�<��<ٽ�<���<���<���<H��<���<q��<��<e��<(��<���<`   `   ��<x��<���<���<l��<j��<h��<���<��<���<u��<���<׽�<���<u��<���<��<���<h��<j��<l��<���<���<x��<`   `   ^��<���<���<��<
��<��<���<��<���<���<G��<V��<���<V��<G��<���<���<��<���<��<
��<��<���<���<`   `   "��< ��<S��<���<7��<r��<P��<���<���<a��<���<��<��<��<���<a��<���<���<P��<r��<7��<���<S��< ��<`   `   ���<(��<���<3��<%��<%��<��<w��<{��<���<*��<b��<��<b��<*��<���<{��<w��<��<%��<%��<3��<���<(��<`   `   ~��<���<���<���<���<���<n��<���<��<%��<���<ػ�<���<ػ�<���<%��<��<���<n��<���<���<���<���<���<`   `   ���<{��<X��<���<I��<���<z��<%��<.��<G��<��<��<��<��<��<G��<.��<%��<z��<���<I��<���<X��<{��<`   `   ���<k��<���<��<8��<���<���<2��<U��<T��<Ǻ�<��<V��<��<Ǻ�<T��<U��<2��<���<���<8��<��<���<k��<`   `   !��<���<��<���<���<���<���<,��<��<L��<���<���<���<���<���<L��<��<,��<���<���<���<���<��<���<`   `   ��<���<���<v��<w��<^��<,��<��<���<Q��<��<ɷ�<
��<ɷ�<��<Q��<���<��<,��<^��<w��<v��<���<���<`   `   =��<��<F��<��<��<5��<��<��<��<f��<��< ��<d��< ��<��<f��<��<��<��<5��<��<��<F��<��<`   `   r��<!��<���<a��<���<��<<��<7��<z��<Ѹ�<G��<���<ƶ�<���<G��<Ѹ�<z��<7��<<��<��<���<a��<���<!��<`   `   ���<���<���<���<U��<��<C��<P��<���<e��<4��<���<���<���<4��<e��<���<P��<C��<��<U��<���<���<���<`   `   /��<��<o��<a��<���<
��<���<��<I��<>��<���<��<���<��<���<>��<I��<��<���<
��<���<a��<o��<��<`   `   ���<���<C��<���<���<��<��<���<���<{��<��<[��<���<[��<��<{��<���<���<��<��<���<���<C��<���<`   `   ¿�<ο�<e��<���<���<���<���<���<��<��<q��<V��<��<V��<q��<��<��<���<���<���<���<���<e��<ο�<`   `   ���<��<���<���<@��<���<7��<3��<���<=��<���<���<���<���<���<=��<���<3��<7��<���<@��<���<���<��<`   `   ��</��<���<ν�<���<\��<���<6��<)��<���<u��<��<ɺ�<��<u��<���<)��<6��<���<\��<���<ν�<���</��<`   `   s��<��<���<���<���<T��<��< ��<F��<B��<i��<��<���<��<i��<B��<F��< ��<��<T��<���<���<���<��<`   `   ��<���<^��<ý�<���<��<Z��<¾�<���<��<I��<-��<'��<-��<I��<��<���<¾�<Z��<��<���<ý�<^��<���<`   `   ���<ܽ�<̽�<��<���<��<���<��<x��<���</��<k��<���<k��</��<���<x��<��<���<��<���<��<̽�<ܽ�<`   `   ���<<��<4��<���<b��<ݿ�<���<4��<&��<���<f��<���<���<���<f��<���<&��<4��<���<ݿ�<b��<���<4��<<��<`   `   L��<׽�<'��<̾�<̿�<���<��<
��<O��<&��<���<��<��<��<���<&��<O��<
��<��<���<̿�<̾�<'��<׽�<`   `   ���<ݽ�<{��<Z��<N��<���<+��<]��<���<���<���<@��<f��<@��<���<���<���<]��<+��<���<N��<Z��<{��<ݽ�<`   `   ��<ٽ�<���<���<���<H��<���<q��<��<e��<(��<���<���<���<(��<e��<��<q��<���<H��<���<���<���<ٽ�<`   `   ׽�<���<u��<���<��<���<h��<j��<l��<���<���<x��<��<x��<���<���<l��<j��<h��<���<��<���<u��<���<`   `   ���<V��<H��<���<���<��<���<��<
��<��<���<���<^��<���<���<��<
��<��<���<��<���<���<H��<V��<`   `   ��<��<���<a��<���<���<P��<r��<7��<���<S��< ��<"��< ��<S��<���<7��<r��<P��<���<���<a��<���<��<`   `   ��<b��<*��<���<{��<w��<��<%��<%��<3��<���<(��<���<(��<���<3��<%��<%��<��<w��<{��<���<*��<b��<`   `   ���<ػ�<���<%��<��<���<n��<���<���<���<���<���<~��<���<���<���<���<���<n��<���<��<%��<���<ػ�<`   `   ��<��<��<G��<.��<%��<z��<���<I��<���<X��<{��<���<{��<X��<���<I��<���<z��<%��<.��<G��<��<��<`   `   V��<��<Ǻ�<T��<U��<2��<���<���<8��<��<���<k��<���<k��<���<��<8��<���<���<2��<U��<T��<Ǻ�<��<`   `   ���<���<���<L��<��<,��<���<���<���<���<��<���<!��<���<��<���<���<���<���<,��<��<L��<���<���<`   `   
��<ɷ�<��<Q��<���<��<,��<^��<w��<v��<���<���<��<���<���<v��<w��<^��<,��<��<���<Q��<��<ɷ�<`   `   d��< ��<��<f��<��<��<��<5��<��<��<F��<��<=��<��<F��<��<��<5��<��<��<��<f��<��< ��<`   `   ƶ�<���<G��<Ѹ�<z��<7��<<��<��<���<a��<���<!��<r��<!��<���<a��<���<��<<��<7��<z��<Ѹ�<G��<���<`   `   ��<��<��<d��<��<.��<���<���<j��<1��<���<���<���<���<���<1��<j��<���<���<.��<��<d��<��<��<`   `   õ�<[��<ݶ�<U��<޹�<���<۽�<���<���<\��<���<���<���<���<���<\��<���<���<۽�<���<޹�<U��<ݶ�<[��<`   `   ���<&��<t��<!��<M��<u��<d��<	��<���<���<���<���<���<���<���<���<���<	��<d��<u��<M��<!��<t��<&��<`   `   ��<6��<���<��<���<���<V��<s��<!��<��<���<��<I��<��<���<��<!��<s��<V��<���<���<��<���<6��<`   `   ��<��<��<���<t��<���<���<I��<���<;��<���<:��<`��<:��<���<;��<���<I��<���<���<t��<���<��<��<`   `   ��<��<��<b��<��<���<���<���<��<c��<���<��<+��<��<���<c��<��<���<���<���<��<b��<��<��<`   `   ���<���<þ�<���<��<��<+��<���<��<���<��<}��<���<}��<��<���<��<���<+��<��<��<���<þ�<���<`   `   ���<���<h��<���<���<���<���<���<��< ��<��<L��<j��<L��<��< ��<��<���<���<���<���<���<h��<���<`   `   ���<j��<E��<���<m��<���<���<j��<���<"��<���<f��<%��<f��<���<"��<���<j��<���<���<m��<���<E��<j��<`   `   ���<���<a��<���<���<���<���<r��<���<���<��<���<H��<���<��<���<���<r��<���<���<���<���<a��<���<`   `   ���<���<���<���<���<���<s��<���<Q��<j��<8��<���<���<���<8��<j��<Q��<���<s��<���<���<���<���<���<`   `   ���<P��<���<s��<���<[��<���<���<��<���<���<��<(��<��<���<���<��<���<���<[��<���<s��<���<P��<`   `   x��<��< ��<���<���<��<���<���<���< ��<���<߿�<���<߿�<���< ��<���<���<���<��<���<���< ��<��<`   `   q��<��<���<���<D��<��<���<���<D��<��<���<���<��<���<���<��<D��<���<���<��<D��<���<���<��<`   `   {��<f��<J��<���<���<���<L��<���<!��<���<���<���<��<���<���<���<!��<���<L��<���<���<���<J��<f��<`   `   ���<]��</��<~��<��<g��<S��<���<���<���<��<���<e��<���<��<���<���<���<S��<g��<��<~��</��<]��<`   `   f��<���<B��<k��<���<��<���<I��<}��<���<��<ý�<���<ý�<��<���<}��<I��<���<��<���<k��<B��<���<`   `   ���<��<��<Q��<���<���<���<���<.��<���<��<Ҽ�<���<Ҽ�<��<���<.��<���<���<���<���<Q��<��<��<`   `   ���<?��<L��<f��<���<���<r��<R��<���<���<Լ�<s��<"��<s��<Լ�<���<���<R��<r��<���<���<f��<L��<?��<`   `   ���<��<���<���< ��<N��<��<��<��<h��<S��<Y��<l��<Y��<S��<h��<��<��<��<N��< ��<���<���<��<`   `   ���<<��<���<���<���<���<���<���<���<��<��<-��<[��<-��<��<��<���<���<���<���<���<���<���<<��<`   `   u��<.��<���<���<���<���<��<��<��<��<?��<ҷ�<n��<ҷ�<?��<��<��<��<��<���<���<���<���<.��<`   `   ��< ��<���<���< ��<7��<���<���<��<��<"��<��<��<��<"��<��<��<���<���<7��< ��<���<���< ��<`   `   ���<���<t��<���<.��<S��<��<P��<��<��<W��<���<õ�<���<W��<��<��<P��<��<S��<.��<���<t��<���<`   `   ���<���<���<1��<j��<���<���<.��<��<d��<��<��<��<��<��<d��<��<.��<���<���<j��<1��<���<���<`   `   ���<���<���<\��<���<���<۽�<���<޹�<U��<ݶ�<[��<õ�<[��<ݶ�<U��<޹�<���<۽�<���<���<\��<���<���<`   `   ���<���<���<���<���<	��<d��<u��<M��<!��<t��<&��<���<&��<t��<!��<M��<u��<d��<	��<���<���<���<���<`   `   I��<��<���<��<!��<s��<V��<���<���<��<���<6��<��<6��<���<��<���<���<V��<s��<!��<��<���<��<`   `   `��<:��<���<;��<���<I��<���<���<t��<���<��<��<��<��<��<���<t��<���<���<I��<���<;��<���<:��<`   `   +��<��<���<c��<��<���<���<���<��<b��<��<��<��<��<��<b��<��<���<���<���<��<c��<���<��<`   `   ���<}��<��<���<��<���<+��<��<��<���<þ�<���<���<���<þ�<���<��<��<+��<���<��<���<��<}��<`   `   j��<L��<��< ��<��<���<���<���<���<���<h��<���<���<���<h��<���<���<���<���<���<��< ��<��<L��<`   `   %��<f��<���<"��<���<j��<���<���<m��<���<E��<j��<���<j��<E��<���<m��<���<���<j��<���<"��<���<f��<`   `   H��<���<��<���<���<r��<���<���<���<���<a��<���<���<���<a��<���<���<���<���<r��<���<���<��<���<`   `   ���<���<8��<j��<Q��<���<s��<���<���<���<���<���<���<���<���<���<���<���<s��<���<Q��<j��<8��<���<`   `   (��<��<���<���<��<���<���<[��<���<s��<���<P��<���<P��<���<s��<���<[��<���<���<��<���<���<��<`   `   ���<߿�<���< ��<���<���<���<��<���<���< ��<��<x��<��< ��<���<���<��<���<���<���< ��<���<߿�<`   `   ��<���<���<��<D��<���<���<��<D��<���<���<��<q��<��<���<���<D��<��<���<���<D��<��<���<���<`   `   ��<���<���<���<!��<���<L��<���<���<���<J��<f��<{��<f��<J��<���<���<���<L��<���<!��<���<���<���<`   `   e��<���<��<���<���<���<S��<g��<��<~��</��<]��<���<]��</��<~��<��<g��<S��<���<���<���<��<���<`   `   ���<ý�<��<���<}��<I��<���<��<���<k��<B��<���<f��<���<B��<k��<���<��<���<I��<}��<���<��<ý�<`   `   ���<Ҽ�<��<���<.��<���<���<���<���<Q��<��<��<���<��<��<Q��<���<���<���<���<.��<���<��<Ҽ�<`   `   "��<s��<Լ�<���<���<R��<r��<���<���<f��<L��<?��<���<?��<L��<f��<���<���<r��<R��<���<���<Լ�<s��<`   `   l��<Y��<S��<h��<��<��<��<N��< ��<���<���<��<���<��<���<���< ��<N��<��<��<��<h��<S��<Y��<`   `   [��<-��<��<��<���<���<���<���<���<���<���<<��<���<<��<���<���<���<���<���<���<���<��<��<-��<`   `   n��<ҷ�<?��<��<��<��<��<���<���<���<���<.��<u��<.��<���<���<���<���<��<��<��<��<?��<ҷ�<`   `   ��<��<"��<��<��<���<���<7��< ��<���<���< ��<��< ��<���<���< ��<7��<���<���<��<��<"��<��<`   `   õ�<���<W��<��<��<P��<��<S��</��<���<t��<���<���<���<t��<���</��<S��<��<P��<��<��<W��<���<`   `   ��<|��<���<���<#��</��<]��<Q��<&��<���<���<t��<���<t��<���<���<&��<Q��<]��</��<#��<���<���<|��<`   `   ���<���<[��<5��<���<.��<���<���<���<R��<��<���<d��<���<��<R��<���<���<���<.��<���<5��<[��<���<`   `   ��<|��<��<a��<>��<���<ҽ�<f��<��<%��<���<���<K��<���<���<%��<��<f��<ҽ�<���<>��<a��<��<|��<`   `   ���<��<��<ݸ�<��<F��<��<���<,��<���<���<r��<���<r��<���<���<,��<���<��<F��<��<ݸ�<��<��<`   `   ��<i��<M��<���<���<4��<F��<)��<���<���<q��<���<U��<���<q��<���<���<)��<F��<4��<���<���<M��<i��<`   `   ���<`��<μ�<���<���<h��<��<���<���<C��<���<��<I��<��<���<C��<���<���<��<h��<���<���<μ�<`��<`   `   ���<���<��<s��<F��<p��<���<���<���<���<?��<Q��<y��<Q��<?��<���<���<���<���<p��<F��<s��<��<���<`   `   ���<���<���<���<��<���<��<���<���<P��<+��<,��<@��<,��<+��<P��<���<���<��<���<��<���<���<���<`   `   ���<���<���<��<��<4��<=��<<��<���<���<V��<"��<��<"��<V��<���<���<<��<=��<4��<��<��<���<���<`   `   8��<��<���<���<u��<D��<���<$��<���<���<���<5��<��<5��<���<���<���<$��<���<D��<u��<���<���<��<`   `   y��<B��<���<��<���<���<���<���<���<y��<A��<b��<`��<b��<A��<y��<���<���<���<���<���<��<���<B��<`   `   ��<���<X��<���<���<1��<<��<x��<��<���<y��<p��<��<p��<y��<���<��<x��<<��<1��<���<���<X��<���<`   `   ���<3��<[��<Q��<��<���<Q��<Z��<���<:��<���<���<���<���<���<:��<���<Z��<Q��<���<��<Q��<[��<3��<`   `   u��<���<���<���<���<)��<���<���<S��<���<l��<���<���<���<l��<���<S��<���<���<)��<���<���<���<���<`   `   ���<���<p��<���<6��<���<���<}��<���<y��<���<���<=��<���<���<y��<���<}��<���<���<6��<���<p��<���<`   `   ���<��<y��<S��<��<y��<���<���<"��<���<v��<ٿ�<��<ٿ�<v��<���<"��<���<���<y��<��<S��<y��<��<`   `   ���<e��<���<.��<1��<���<���<���<4��<���<���<־�<f��<־�<���<���<4��<���<���<���<1��<.��<���<e��<`   `   ]��<A��<���<���<q��<���<��<���<-��<���<��<L��<Y��<L��<��<���<-��<���<��<���<q��<���<���<A��<`   `   R��<���<��<g��<���<��<���<���<���<h��<���<���<M��<���<���<h��<���<���<���<��<���<g��<��<���<`   `   ���<���<,��<���<8��<H��<���<���<���<z��<��<��<��<��<��<z��<���<���<���<H��<8��<���<,��<���<`   `   :��<���<C��<���<!��<��<���<���<ӿ�<e��<3��<k��<C��<k��<3��<e��<ӿ�<���<���<��<!��<���<C��<���<`   `   $��<���<s��<���<���<���<���<���<D��<���<I��<۶�<ĵ�<۶�<I��<���<D��<���<���<���<���<���<s��<���<`   `   t��<���<j��<���<���<c��<���<���<_��<��<���<���<���<���<���<��<_��<���<���<c��<���<���<j��<���<`   `   ���<	��<���<,��<q��<7��<���<��<���<��<���<޴�<?��<޴�<���<��<���<��<���<7��<q��<,��<���<	��<`   `   ���<t��<���<���<&��<Q��<]��</��<#��<���<���<|��<��<|��<���<���<#��</��<]��<Q��<&��<���<���<t��<`   `   d��<���<��<R��<���<���<���<.��<���<5��<[��<���<���<���<[��<5��<���<.��<���<���<���<R��<��<���<`   `   K��<���<���<%��<��<f��<ҽ�<���<>��<a��<��<|��<��<|��<��<a��<>��<���<ҽ�<f��<��<%��<���<���<`   `   ���<r��<���<���<,��<���<��<F��<��<ݸ�<��<��<���<��<��<ݸ�<��<F��<��<���<,��<���<���<r��<`   `   U��<���<q��<���<���<)��<F��<4��<���<���<M��<i��<��<i��<M��<���<���<4��<F��<)��<���<���<q��<���<`   `   I��<��<���<C��<���<���<��<h��<���<���<μ�<`��<���<`��<μ�<���<���<h��<��<���<���<C��<���<��<`   `   x��<Q��<?��<���<���<���<���<p��<F��<s��<��<���<���<���<��<s��<F��<p��<���<���<���<���<?��<Q��<`   `   @��<,��<+��<P��<���<���<��<���<��<���<���<���<���<���<���<���<��<���<��<���<���<P��<+��<,��<`   `   ��<"��<V��<���<���<<��<=��<4��<��<��<���<���<���<���<���<��<��<4��<=��<<��<���<���<V��<"��<`   `   ��<5��<���<���<���<$��<���<D��<u��<���<���<��<8��<��<���<���<u��<D��<���<$��<���<���<���<5��<`   `   `��<b��<A��<y��<���<���<���<���<���<��<���<B��<y��<B��<���<��<���<���<���<���<���<y��<A��<b��<`   `   ��<p��<y��<���<��<x��<<��<1��<���<���<X��<���<��<���<X��<���<���<1��<<��<x��<��<���<y��<p��<`   `   ���<���<���<:��<���<Z��<Q��<���<��<Q��<[��<3��<���<3��<[��<Q��<��<���<Q��<Z��<���<:��<���<���<`   `   ���<���<l��<���<S��<���<���<)��<���<���<���<���<u��<���<���<���<���<)��<���<���<S��<���<l��<���<`   `   =��<���<���<y��<���<}��<���<���<6��<���<p��<���<���<���<p��<���<6��<���<���<}��<���<y��<���<���<`   `   ��<ٿ�<v��<���<"��<���<���<y��<��<S��<y��<��<���<��<y��<S��<��<y��<���<���<"��<���<v��<ٿ�<`   `   f��<־�<���<���<4��<���<���<���<1��<.��<���<e��<���<e��<���<.��<1��<���<���<���<4��<���<���<־�<`   `   Y��<L��<��<���<-��<���<��<���<q��<���<���<A��<]��<A��<���<���<q��<���<��<���<-��<���<��<L��<`   `   M��<���<���<h��<���<���<���<��<���<g��<��<���<R��<���<��<g��<���<��<���<���<���<h��<���<���<`   `   ��<��<��<z��<���<���<���<H��<8��<���<,��<���<���<���<,��<���<8��<H��<���<���<���<z��<��<��<`   `   C��<k��<3��<e��<Կ�<���<���<��<!��<���<C��<���<:��<���<C��<���<!��<��<���<���<Կ�<e��<3��<k��<`   `   ĵ�<۶�<I��<���<D��<���<���<���<���<���<s��<���<$��<���<s��<���<���<���<���<���<D��<���<I��<۶�<`   `   ���<���<���<��<_��<���<���<c��<���<���<j��<���<t��<���<j��<���<���<c��<���<���<_��<��<���<���<`   `   ?��<޴�<���<��<���<��<���<7��<q��<,��<���<	��<���<	��<���<,��<q��<7��<���<��<���<��<���<޴�<`   `   ���<���<���<��<E��<`��<~��<��<���<,��<���<���<n��<���<���<,��<���<��<~��<`��<E��<��<���<���<`   `   ���<��<C��<)��<ڷ�<b��<þ�<���<7��<5��<B��<���<���<���<B��<5��<7��<���<þ�<b��<ڷ�<)��<C��<��<`   `   ��<���<g��<յ�<e��<M��<��<p��<Y��<���<���<���<��<���<���<���<Y��<p��<��<M��<e��<յ�<g��<���<`   `   ��<���<���<��<���<z��<���<���<���<���<E��<��<8��<��<E��<���<���<���<���<z��<���<��<���<���<`   `   ���<���<?��<���<P��<Z��<0��<r��<���<���<^��<���<���<���<^��<���<���<r��<0��<Z��<P��<���<?��<���<`   `   ̻�<��<*��<���<���<z��<տ�<���<���<���<7��<���<���<���<7��<���<���<���<տ�<z��<���<���<*��<��<`   `   _��<���<���<���<���<d��<���<���<B��<J��<4��<���<}��<���<4��<J��<B��<���<���<d��<���<���<���<���<`   `   ���<��<���<B��<��<���<%��<8��<5��<���<+��<7��<���<7��<+��<���<5��<8��<%��<���<��<B��<���<��<`   `   ���<���<���<���<��<��<��<���<���<���<���<+��<���<+��<���<���<���<���<��<��<��<���<���<���<`   `   @��<��<��<���<N��<d��<���<���<���<b��<-��<8��<��<8��<-��<b��<���<���<���<d��<N��<���<��<��<`   `   ��<`��<b��<���<���<'��<Y��<���<K��<9��<���<���<i��<���<���<9��<K��<���<Y��<'��<���<���<b��<`��<`   `   m��<|��<��<��<|��<���<`��<
��<���<��<8��<���<<��<���<8��<��<���<
��<`��<���<|��<��<��<|��<`   `   ���<	��<x��<���<���<���<q��<���<���<���<���<��<J��<��<���<���<���<���<q��<���<���<���<x��<	��<`   `   ��<���<1��<@��<��<E��<���<���<i��<<��<.��<���<+��<���<.��<<��<i��<���<���<E��<��<@��<1��<���<`   `   ��<���<���<R��<���<���<��<2��<���< ��<���<���<g��<���<���< ��<���<2��<��<���<���<R��<���<���<`   `   ���<H��<��<���<K��<L��<a��<��<���<��<���<��<k��<��<���<��<���<��<a��<L��<K��<���<��<H��<`   `   (��<���<y��<��<x��<D��<���<=��<���<���<t��<"��<M��<"��<t��<���<���<=��<���<D��<x��<��<y��<���<`   `   ���<$��<���<.��<l��<��<w��<���<���<���<j��<��<)��<��<j��<���<���<���<w��<��<l��<.��<���<$��<`   `   M��<���<���<���<���<@��<���<���<o��<|��<-��<b��<���<b��<-��<|��<o��<���<���<@��<���<���<���<���<`   `   s��<���<���</��<���<��<r��<���<��<;��<̺�<���<(��<���<̺�<;��<��<���<r��<��<���</��<���<���<`   `   i��<���<Y��<���<*��<��<���<���<���<��<T��<k��<���<k��<T��<��<���<���<���<��<*��<���<Y��<���<`   `   ��<���<���<&��<���<��<���<���<��<ҹ�<E��<���<@��<���<E��<ҹ�<��<���<���<��<���<&��<���<���<`   `   ���<y��<���<���<r��<���<���<���<���<��<д�<���<��<���<д�<��<���<���<���<���<r��<���<���<y��<`   `   ��<z��<���<���<���<���<���<I��<չ�<h��<U��<��<���<��<U��<h��<չ�<I��<���<���<���<���<���<z��<`   `   n��<���<���<,��<���<��<~��<`��<E��<��<���<���<���<���<���<��<E��<`��<~��<��<���<,��<���<���<`   `   ���<���<B��<5��<7��<���<þ�<a��<ڷ�<)��<C��<��<���<��<C��<)��<ڷ�<a��<þ�<���<7��<5��<B��<���<`   `   ��<���<���<���<Y��<p��<��<M��<e��<յ�<f��<���<��<���<f��<յ�<e��<M��<��<p��<Y��<���<���<���<`   `   8��<��<E��<���<���<���<���<z��<���<��<���<���<��<���<���<��<���<z��<���<���<���<���<E��<��<`   `   ���<���<^��<���<���<r��<0��<Z��<P��<���<?��<���<���<���<?��<���<P��<Z��<0��<r��<���<���<^��<���<`   `   ���<���<7��<���<���<���<տ�<z��<���<���<*��<��<̻�<��<*��<���<���<z��<տ�<���<���<���<7��<���<`   `   }��<���<4��<J��<B��<���<���<d��<���<���<���<���<_��<���<���<���<���<d��<���<���<B��<J��<4��<���<`   `   ���<7��<+��<���<5��<8��<%��<���<��<B��<���<��<���<��<���<B��<��<���<%��<8��<5��<���<+��<7��<`   `   ���<+��<���<���<���<���<��<��<��<���<���<���<���<���<���<���<��<��<��<���<���<���<���<+��<`   `   ��<8��<-��<b��<���<���<���<d��<N��<���<��<��<@��<��<��<���<N��<d��<���<���<���<b��<-��<8��<`   `   i��<���<���<9��<K��<���<Y��<'��<���<���<b��<`��<��<`��<b��<���<���<'��<Y��<���<K��<9��<���<���<`   `   <��<���<8��<��<���<
��<`��<���<|��<��<��<|��<m��<|��<��<��<|��<���<`��<
��<���<��<8��<���<`   `   J��<��<���<���<���<���<q��<���<���<���<x��<	��<���<	��<x��<���<���<���<q��<���<���<���<���<��<`   `   +��<���<.��<<��<i��<���<���<E��<��<@��<1��<���<��<���<1��<@��<��<E��<���<���<i��<<��<.��<���<`   `   g��<���<���< ��<���<2��<��<���<���<R��<���<���<��<���<���<R��<���<���<��<2��<���< ��<���<���<`   `   k��<��<���<��<���<��<a��<L��<K��<���<��<H��<���<H��<��<���<K��<L��<a��<��<���<��<���<��<`   `   M��<"��<t��<���<���<=��<���<D��<x��<��<y��<���<(��<���<y��<��<x��<D��<���<=��<���<���<t��<"��<`   `   )��<��<j��<���<���<���<w��<��<l��<.��<���<$��<���<$��<���<.��<l��<��<w��<���<���<���<j��<��<`   `   ���<b��<-��<|��<o��<���<���<A��<���<���<���<���<M��<���<���<���<���<A��<���<���<o��<|��<-��<b��<`   `   (��<���<̺�<;��<��<���<r��<��<���</��<���<���<s��<���<���</��<���<��<r��<���<��<;��<̺�<���<`   `   ���<k��<T��<��<���<���<���<��<*��<���<Y��<���<i��<���<Y��<���<*��<��<���<���<���<��<T��<k��<`   `   @��<���<E��<ҹ�<��<���<���<��<���<&��<���<���<��<���<���<&��<���<��<���<���<��<ҹ�<E��<���<`   `   ��<���<Ѵ�<��<���<���<���<���<r��<���<���<y��<���<y��<���<���<r��<���<���<���<���<��<Ѵ�<���<`   `   ���<��<U��<h��<չ�<J��<���<���<���<���<���<z��<��<z��<���<���<���<���<���<J��<չ�<h��<U��<��<`   `   h��<���<���<��<��<��<���<���<��<���<"��<���<���<���<"��<���<��<���<���<��<��<��<���<���<`   `   ���<��<ɭ�<���<��<{��<���<V��<��<6��<.��<~��<���<~��<.��<6��<��<V��<���<{��<��<���<ɭ�<��<`   `   P��<���<$��<���<��<��<���<��<!��<���<���<���<���<���<���<���<!��<��<���<��<��<���<$��<���<`   `   ���<���<ӱ�<��<W��<U��<��<���<@��<���<���<s��<���<s��<���<���<@��<���<��<U��<W��<��<ӱ�<���<`   `   Q��<״�<���<W��<0��<:��<½�<���<��<"��<[��<`��<���<`��<[��<"��<��<���<½�<:��<0��<W��<���<״�<`   `   Ϲ�<w��<(��<���<��<��<\��<w��<���<��<���<n��<���<n��<���<��<���<w��<\��<��<��<���<(��<w��<`   `   ���<���<���<���<@��<P��<���<��<k��<���<M��<y��<H��<y��<M��<���<k��<��<���<P��<@��<���<���<���<`   `   ���<���<N��<��<e��<v��<%��<���<���<m��<J��<���<���<���<J��<m��<���<���<%��<v��<e��<��<N��<���<`   `   '��<��<w��<���<G��<e��<���<��<J��<5��<t��<���<���<���<t��<5��<J��<��<���<e��<G��<���<w��<��<`   `   ���<���<���<I��<��<n��<q��<���<���<{��<���<���<���<���<���<{��<���<���<q��<n��<��<I��<���<���<`   `   ���<;��<���<���<z��<|��<���<��<��<���<���<���<��<���<���<���<��<��<���<|��<z��<���<���<;��<`   `   ���<��<[��<���<���<���<���<R��<���<O��<<��<���<N��<���<<��<O��<���<R��<���<���<���<���<[��<��<`   `   ���<0��<-��<���<���<R��<1��<���<���<��<s��<���<��<���<s��<��<���<���<1��<R��<���<���<-��<0��<`   `   ��<0��<���<���<}��<q��<���<��<���<��<���<>��<��<>��<���<��<���<��<���<q��<}��<���<���<0��<`   `   v��<w��<5��<���<���<���<���<���<���<���<��<I��<���<I��<��<���<���<���<���<���<���<���<5��<w��<`   `   ���<���<1��<���< ��<_��<���<���<���<���<H��<���<��<���<H��<���<���<���<���<_��< ��<���<1��<���<`   `   ���<w��<���<Y��<*��<���<���<&��<;��<��<<��<���<��<���<<��<��<;��<&��<���<���<*��<Y��<���<w��<`   `   ���<���<���<��<���<���<���<��<��<���<J��<K��<��<K��<J��<���<��<��<���<���<���<��<���<���<`   `   \��<���<���<���<\��<��<9��<C��<+��<���<9��<!��<·�<!��<9��<���<+��<C��<9��<��<\��<���<���<���<`   `   $��<V��<a��<M��<���<���<���<(��<���<��<���<��<Ӵ�<��<���<��<���<(��<���<���<���<M��<a��<V��<`   `   ���<���<���<��<��<���<��<���<���<���<��<���<ر�<���<��<���<���<���<��<���<��<��<���<���<`   `   ���<���<��<~��<���<���<&��<���<��<@��<���<���<ڮ�<���<���<@��<��<���<&��<���<���<~��<��<���<`   `   R��<a��<���<R��<���<.��<5��<���<ڹ�<C��<u��<���<���<���<u��<C��<ڹ�<���<5��<.��<���<R��<���<a��<`   `   ��<���<���<<��<N��<<��<���<Խ�<���<D��<Ԯ�<9��<t��<9��<Ԯ�<D��<���<Խ�<���<<��<N��<<��<���<���<`   `   ���<���<!��<���<��<���<���<��<��<��<���<���<h��<���<���<��<��<��<���<���<��<���<!��<���<`   `   ���<~��<.��<6��<��<V��<���<{��<��<���<ɭ�<��<���<��<ɭ�<���<��<{��<���<V��<��<6��<.��<~��<`   `   ���<���<���<���<!��<��<���<��<��<���<$��<���<P��<���<$��<���<��<��<���<��<!��<���<���<���<`   `   ���<s��<���<���<@��<���<��<U��<W��<��<ӱ�<���<���<���<ӱ�<��<W��<U��<��<���<@��<���<���<s��<`   `   ���<`��<[��<"��<��<���<½�<:��<0��<W��<���<ִ�<Q��<ִ�<���<W��<0��<:��<½�<���<��<"��<[��<`��<`   `   ���<n��<���<��<���<w��<\��<��<��<���<(��<w��<Ϲ�<w��<(��<���<��<��<\��<w��<���<��<���<n��<`   `   H��<y��<M��<���<k��<��<���<P��<@��<���<���<���<���<���<���<���<@��<P��<���<��<k��<���<M��<y��<`   `   ���<���<J��<m��<���<���<%��<v��<e��<��<N��<���<���<���<N��<��<e��<v��<%��<���<���<m��<J��<���<`   `   ���<���<t��<5��<J��<��<���<e��<G��<���<w��<��<'��<��<w��<���<G��<e��<���<��<J��<5��<t��<���<`   `   ���<���<���<{��<���<���<q��<n��<��<I��<���<���<���<���<���<I��<��<n��<q��<���<���<{��<���<���<`   `   ��<���<���<���<��<��<���<|��<z��<���<���<;��<���<;��<���<���<z��<|��<���<��<��<���<���<���<`   `   N��<���<<��<O��<���<R��<���<���<���<���<[��<��<���<��<[��<���<���<���<���<R��<���<O��<<��<���<`   `   ��<���<s��<��<���<���<1��<R��<���<���<-��<0��<���<0��<-��<���<���<R��<1��<���<���<��<s��<���<`   `   ��<>��<���<��<���<��<���<q��<}��<���<���<0��<��<0��<���<���<}��<q��<���<��<���<��<���<>��<`   `   ���<I��<��<���<���<���<���<���<���<���<5��<w��<v��<w��<5��<���<���<���<���<���<���<���<��<I��<`   `   ��<���<H��<���<���<���<���<_��< ��<���<1��<���<���<���<1��<���< ��<_��<���<���<���<���<H��<���<`   `   ��<���<<��<��<;��<&��<���<���<*��<Y��<���<w��<���<w��<���<Y��<*��<���<���<&��<;��<��<<��<���<`   `   ��<K��<J��<���<��<��<���<���<���<��<���<���<���<���<���<��<���<���<���<��<��<���<J��<K��<`   `   ·�<!��<9��<���<+��<C��<9��<��<\��<���<���<���<\��<���<���<���<\��<��<9��<C��<+��<���<9��<!��<`   `   Ӵ�<��<���<��<���<(��<���<���<���<M��<a��<V��<$��<V��<a��<M��<���<���<���<(��<���<��<���<��<`   `   ر�<���<��<���<���<���<��<���<��<��<���<���<���<���<���<��<��<���<��<���<���<���<��<���<`   `   ڮ�<���<���<@��<��<���<&��<���<���<~��<��<���<���<���<��<~��<���<���<&��<���<��<@��<���<���<`   `   ���<���<u��<C��<ڹ�<���<5��<.��<���<R��<���<a��<R��<a��<���<R��<���<.��<5��<���<ڹ�<C��<u��<���<`   `   t��<9��<ծ�<D��<���<Խ�<���<<��<N��<<��<���<���<��<���<���<<��<N��<<��<���<Խ�<���<D��<ծ�<9��<`   `   ���<��<\��<"��<=��<��<���<m��<���<��<r��<���<���<���<r��<��<���<m��<���<��<=��<"��<\��<��<`   `   ���<��<���<���<=��<���<��<���<���<_��<v��<.��<���<.��<v��<_��<���<���<��<���<=��<���<���<��<`   `   k��<X��<6��<��<M��<��<��<���<��<a��<��<~��<���<~��<��<a��<��<���<��<��<M��<��<6��<X��<`   `   ���<A��<%��<��<���<F��<���<ʾ�<U��<���<���<j��<���<j��<���<���<U��<ʾ�<���<F��<���<��<%��<A��<`   `   ���<ݯ�<J��<���<0��<���<���<���<���<���<N��<L��<���<L��<N��<���<���<���<���<���<0��<���<J��<ݯ�<`   `   -��<��<���<���<��<���<���<¿�<���<��<��<���<U��<���<��<��<���<¿�<���<���<��<���<���<��<`   `   ���<M��<���<,��<���<���<B��<(��<��<���<���<U��<q��<U��<���<���<��<(��<B��<���<���<,��<���<M��<`   `   ���<���<���<A��<H��<���<���<��<)��<b��<���<h��<p��<h��<���<b��<)��<��<���<���<H��<A��<���<���<`   `   ���<2��<c��<���<���<��<���<j��<a��<���<E��<l��<���<l��<E��<���<a��<j��<���<��<���<���<c��<2��<`   `   ��<���<���<���<���<���<3��<���<M��<���<~��<���<���<���<~��<���<M��<���<3��<���<���<���<���<���<`   `   5��<���<[��<U��<}��<���<<��<���<��<���<���<x��<^��<x��<���<���<��<���<<��<���<}��<U��<[��<���<`   `   T��<��<m��<���<���<���<���<��<���<���< ��<���<���<���< ��<���<���<��<���<���<���<���<m��<��<`   `   ���<���<��<���<��<���<:��<���<���<��<n��<���<	��<���<n��<��<���<���<:��<���<��<���<��<���<`   `   �<t��<b��<I��<q��<���<6��< ��<���<@��<\��<��<{��<��<\��<@��<���< ��<6��<���<q��<I��<b��<t��<`   `   c�<��<p�<���<���<&��<���<���< ��<���<h��<F��<���<F��<h��<���< ��<���<���<&��<���<���<p�<��<`   `   &	�<��<�<���<���<@��<l��<���<��<e��<q��<ٿ�<��<ٿ�<q��<e��<��<���<l��<@��<���<���<�<��<`   `   
�<��<s�<���<���<���<f��<F��<���<���<���<���<���<���<���<���<���<F��<f��<���<���<���<s�<��<`   `   ��<��<��<���<l��<���<���<���<���<���<���<���<g��<���<���<���<���<���<���<���<l��<���<��<��<`   `   ��<Z�<h �<���<)��<���<���<@��<���<��<n��<C��</��<C��<n��<��<���<@��<���<���<)��<���<h �<Z�<`   `   ��<���<z��<���<���<��<V��<���<���<���<@��<L��<.��<L��<@��<���<���<���<V��<��<���<���<z��<���<`   `   ���<���<���<���<r��<���<c��<��<$��<���<C��<���< ��<���<C��<���<$��<��<c��<���<r��<���<���<���<`   `   ���<���<'��< ��< ��<���<��<M��<[��<��<*��<���<��<���<*��<��<[��<M��<��<���< ��< ��<'��<���<`   `   ���<���<��<���<\��< ��<���<#��<���<]��<���<p��<P��<p��<���<]��<���<#��<���< ��<\��<���<��<���<`   `   u��<A��<}��<V��<Z��<���<���<��<6��<��<T��<���<��<���<T��<��<6��<��<���<���<Z��<V��<}��<A��<`   `   ���<���<r��<��<���<m��<���<��<=��<"��<\��<��<���<��<\��<"��<=��<��<���<m��<���<��<r��<���<`   `   ���<.��<v��<_��<���<���<��<���<=��<���<���<��<���<��<���<���<=��<���<��<���<���<_��<v��<.��<`   `   ���<~��<��<a��<��<���<��<��<M��<��<6��<X��<k��<X��<6��<��<M��<��<��<���<��<a��<��<~��<`   `   ���<j��<���<���<U��<ʾ�<���<F��<���<��<%��<A��<���<A��<%��<��<���<F��<���<ʾ�<U��<���<���<j��<`   `   ���<L��<N��<���<���<���<���<���<0��<���<J��<ݯ�<���<ݯ�<J��<���<0��<���<���<���<���<���<N��<L��<`   `   U��<���<��<��<���<¿�<���<���<��<���<���<��<-��<��<���<���<��<���<���<¿�<���<��<��<���<`   `   q��<U��<���<���<��<'��<B��<���<���<,��<���<M��<���<M��<���<,��<���<���<B��<'��<��<���<���<U��<`   `   p��<h��<���<b��<)��<��<���<���<H��<@��<���<���<���<���<���<@��<H��<���<���<��<)��<b��<���<h��<`   `   ���<l��<E��<���<a��<j��<���<��<���<���<c��<2��<���<2��<c��<���<���<��<���<j��<a��<���<E��<l��<`   `   ���<���<~��<���<M��<���<3��<���<���<���<���<���<��<���<���<���<���<���<3��<���<M��<���<~��<���<`   `   ^��<x��<���<���<��<���<<��<���<}��<U��<[��<���<5��<���<[��<U��<}��<���<<��<���<��<���<���<x��<`   `   ���<���< ��<���<���<��<���<���<���<���<m��<��<T��<��<m��<���<���<���<���<��<���<���< ��<���<`   `   	��<���<n��<��<���<���<:��<���<��<���<��<���<���<���<��<���<��<���<:��<���<���<��<n��<���<`   `   {��<��<\��<@��<���< ��<6��<���<q��<I��<b��<t��<�<t��<b��<I��<q��<���<6��< ��<���<@��<\��<��<`   `   ���<F��<h��<���< ��<���<���<&��<���<���<q�<��<c�<��<q�<���<���<&��<���<���< ��<���<h��<F��<`   `   ��<ٿ�<q��<e��<��<���<l��<@��<���<���<�<��<&	�<��<�<���<���<@��<l��<���<��<e��<q��<ٿ�<`   `   ���<���<���<���<���<F��<f��<���<���<���<s�<��<
�<��<s�<���<���<���<f��<F��<���<���<���<���<`   `   g��<���<���<���<���<���<���<���<l��<���<��<��<��<��<��<���<l��<���<���<���<���<���<���<���<`   `   /��<C��<n��<��<���<@��<���<���<)��<���<h �<Z�<��<Z�<h �<���<)��<���<���<@��<���<��<n��<C��<`   `   .��<L��<@��<���<���<���<W��<��<���<���<z��<���<��<���<z��<���<���<��<W��<���<���<���<@��<L��<`   `    ��<���<C��<���<$��<��<c��<���<r��<���<���<���<���<���<���<���<r��<���<c��<��<$��<���<C��<���<`   `   ��<���<*��<��<\��<M��<��<���< ��< ��<'��<���<���<���<'��< ��< ��<���<��<M��<\��<��<*��<���<`   `   P��<p��<���<]��<���<#��<���< ��<\��<���<��<���<���<���<��<���<\��< ��<���<#��<���<]��<���<p��<`   `   ��<���<T��<��<6��<��<���<���<Z��<V��<}��<A��<u��<A��<}��<V��<Z��<���<���<��<6��<��<T��<���<`   `   ���<0��<��<��<4��<_��<r��<���<p��<���<~��<w��<7��<w��<~��<���<p��<���<r��<_��<4��<��<��<0��<`   `   ��<L��<\��<}��<ҧ�<��<B��<���<��<C��<���<I��<$��<I��<���<C��<��<���<B��<��<ҧ�<}��<\��<L��<`   `   ڙ�<1��<ѝ�<W��<���<���<Ŷ�<Ҿ�<���<���<���<-��<���<-��<���<���<���<Ҿ�<Ŷ�<���<���<W��<ѝ�<1��<`   `   ���<u��<~��<0��<��<���<?��<���<���<}��<���<���<���<���<���<}��<���<���<?��<���<��<0��<~��<u��<`   `   ӧ�<'��<f��<)��<���<���<���<6��<ٿ�<$��<y��<���<���<���<y��<$��<ٿ�<6��<���<���<���<)��<f��<'��<`   `   ���<б�<���<S��<��</��<���<m��<���<���<���<���<���<���<���<���<���<m��<���</��<��<S��<���<б�<`   `   ���<6��<���<���<2��<���<���<���<���<���<$��<l��<4��<l��<$��<���<���<���<���<���<2��<���<���<6��<`   `   ��<���<���<��<���<���<B��<���<��<q��<���<���<#��<���<���<q��<��<���<B��<���<���<��<���<���<`   `   ��<���<���<���<��<��<��<H��<���<Q��<w��<o��<���<o��<w��<Q��<���<H��<��<��<��<���<���<���<`   `   ��<Z��<���<��<���<��<n��<���<��<���<���<���<O��<���<���<���<��<���<n��<��<���<��<���<Z��<`   `   ���<��<t��<���<v��<���<K��<���<���<���<���<���<
��<���<���<���<���<���<K��<���<v��<���<t��<��<`   `   � �< �<f��<]��<���<��<��<"��<[��<���<M��<��<=��<��<M��<���<[��<"��<��<��<���<]��<f��< �<`   `   #�<8�<�<� �<��<*��<���<��<���<9��<���<���<���<���<���<9��<���<��<���<*��<��<� �<�<8�<`   `   R�<��<��<	�<���<���<{��<s��<{��<���<K��<���<���<���<K��<���<{��<s��<{��<���<���<	�<��<��<`   `   #�<s�<��<��<��<��<��<���<���<'��<���<��<Ͼ�<��<���<'��<���<���<��<��<��<��<��<s�<`   `    �<��<H�<V�<��<y��<���<���<{��<P��<���<���<��<���<���<P��<{��<���<���<y��<��<V�<H�<��<`   `   !�<��<\�<��<�<���<���<���<��<m��<8��<���<���<���<8��<m��<��<���<���<���<�<��<\�<��<`   `   ' �<B�<��<V�<��<8��<)��<[��<��<���<4��<��<��<��<4��<���<��<[��<)��<8��<��<V�<��<B�<`   `   T�<�<��<�<4 �<���<b��<l��<��<ƽ�<��<���<"��<���<��<ƽ�<��<l��<b��<���<4 �<�<��<�<`   `   ��<��<��<��<��<���<u��<u��<h��<A��<p��<ߩ�<-��<ߩ�<p��<A��<h��<u��<u��<���<��<��<��<��<`   `   -�<V�<��<��<���<���<���<���<��<��<c��<#��<=��<#��<c��<��<��<���<���<���<���<��<��<V�<`   `   ��<��<M��<��<7��<���<���<���<��<e��<9��<!��<��<!��<9��<e��<��<���<���<���<7��<��<M��<��<`   `   ��<��<���<P��<��</��<���<̼�<l��<���<ş�<���<���<���<ş�<���<l��<̼�<���</��<��<P��<���<��<`   `   ���<s��<3��<1��<���<z��<!��<���<���<���<x��<��<��<��<x��<���<���<���<!��<z��<���<1��<3��<s��<`   `   7��<w��<~��<���<p��<���<r��<_��<4��<��<��<0��<���<0��<��<��<4��<_��<r��<���<p��<���<~��<w��<`   `   $��<I��<���<C��<��<���<B��<��<ѧ�<}��<\��<L��<��<L��<\��<}��<ѧ�<��<B��<���<��<C��<���<I��<`   `   ���<-��<���<���<���<Ҿ�<Ŷ�<���<���<W��<ѝ�<0��<ڙ�<0��<ѝ�<W��<���<���<Ŷ�<Ҿ�<���<���<���<-��<`   `   ���<���<���<}��<���<���<?��<���<��<0��<~��<u��<���<u��<~��<0��<��<���<?��<���<���<}��<���<���<`   `   ���<���<y��<$��<ٿ�<6��<���<���<���<)��<e��<&��<ӧ�<&��<e��<)��<���<���<���<6��<ٿ�<$��<y��<���<`   `   ���<���<���<���<���<m��<���</��<��<S��<���<б�<���<б�<���<S��<��</��<���<m��<���<���<���<���<`   `   4��<l��<$��<���<���<���<���<���<2��<���<���<6��<���<6��<���<���<2��<���<���<���<���<���<$��<l��<`   `   #��<���<���<q��<��<���<B��<���<���<��<���<���<��<���<���<��<���<���<B��<���<��<q��<���<���<`   `   ���<o��<w��<Q��<���<H��<��<��<��<���<���<���<��<���<���<���<��<��<��<H��<���<Q��<w��<o��<`   `   O��<���<���<���<��<���<n��<��<���<��<���<Z��<��<Z��<���<��<���<��<n��<���<��<���<���<���<`   `   
��<���<���<���<���<���<K��<���<v��<���<t��<��<���<��<t��<���<v��<���<K��<���<���<���<���<���<`   `   =��<��<M��<���<[��<"��<��<��<���<]��<f��< �<� �< �<f��<]��<���<��<��<"��<[��<���<M��<��<`   `   ���<���<���<9��<���<��<���<*��<��<� �<�<8�<#�<8�<�<� �<��<*��<���<��<���<9��<���<���<`   `   ���<���<K��<���<{��<s��<{��<���<���<	�<��<��<S�<��<��<	�<���<���<{��<s��<{��<���<K��<���<`   `   Ͼ�<��<���<'��<���<���<��<��<��<��<��<s�<#�<s�<��<��<��<��<��<���<���<'��<���<��<`   `   ��<���<���<P��<{��<���<���<y��<��<V�<H�<��< �<��<H�<V�<��<y��<���<���<{��<P��<���<���<`   `   ���<���<8��<m��<��<���<���<���<�<��<\�<��<!�<��<\�<��<�<���<���<���<��<m��<8��<���<`   `   ��<��<4��<���<��<[��<)��<8��<��<V�<��<B�<' �<B�<��<V�<��<8��<)��<[��<��<���<4��<��<`   `   "��<���<��<ƽ�<��<m��<b��<���<4 �<�<��<�<T�<�<��<�<4 �<���<b��<m��<��<ƽ�<��<���<`   `   -��<ߩ�<p��<A��<h��<u��<u��<���<��<��<��<��<��<��<��<��<��<���<u��<u��<h��<A��<p��<ߩ�<`   `   =��<$��<c��<��<��<���<���<���<���<��<��<V�<.�<V�<��<��<���<���<���<���<��<��<c��<$��<`   `   ��<!��<:��<e��<��<���<���<���<7��<��<M��<��<��<��<M��<��<7��<���<���<���<��<e��<:��<!��<`   `   ���<���<ş�<���<l��<̼�<���</��<��<P��<���<��<��<��<���<P��<��</��<���<̼�<l��<���<ş�<���<`   `   ��<��<x��<���<���<���<!��<z��<���<1��<3��<s��<���<s��<3��<1��<���<z��<!��<���<���<���<x��<��<`   `   ��<���<��<���<w��<���<��<���<���<|��<���< ��<���< ��<���<|��<���<���<��<���<w��<���<��<���<`   `   D��<���<_��<3��<h��<��<ӳ�<'��<o��<H��<F��<���<���<���<F��<H��<o��<'��<ӳ�<��<h��<3��<_��<���<`   `   ǉ�<��<��<z��<��<���<���<���<���<���<?��<���<���<���<?��<���<���<���<���<���<��<z��<��<��<`   `   E��<v��<v��</��<���<���<��<��<���<y��<H��<+��<���<+��<H��<y��<���<��<��<���<���</��<v��<v��<`   `   |��<���<���<.��<���<ʫ�<���<e��<��<���<6��<���<���<���<6��<���<��<e��<���<ʫ�<���<.��<���<���<`   `   ���<���<��<���<���<a��< ��<"��<���<i��<5��<���<.��<���<5��<i��<���<"��< ��<a��<���<���<��<���<`   `   ���<5��<>��<~��<0��<Ϻ�<U��<#��<H��<(��<U��<���<)��<���<U��<(��<H��<#��<U��<Ϻ�<0��<~��<>��<5��<`   `   t��<U��<@��<T��<p��<_��<��<���<W��<��<'��<��<���<��<'��<��<W��<���<��<_��<p��<T��<@��<U��<`   `   @��<���<���<T��<e��<��<>��<���<���<5��<9��<���<Խ�<���<9��<5��<���<���<>��<��<e��<T��<���<���<`   `   ���<��<���<L��<���<.��<��<���<���<���<���<���<���<���<���<���<���<���<��<.��<���<L��<���<��<`   `   �<��<Q��<t��<#��<���<���<���<��<T��<Q��</��<y��</��<Q��<T��<��<���<���<���<"��<t��<Q��<��<`   `   �<u�<J�<�<e��<\��<6��<N��<���<���<���<���<���<���<���<���<���<N��<6��<\��<e��<�<J�<u�<`   `   V#�<�!�<��<y�<�	�<|��<_��<���<y��<9��<���<���<p��<���<���<9��<y��<���<_��<|��<�	�<y�<��<�!�<`   `   �/�<U.�<7(�<��<�<�<0��<���<���<J��<���<��<O��<��<���<J��<���<���<0��<�<�<��<7(�<U.�<`   `   �8�<v7�<`0�<�%�<7�<�	�<���<c��<@��<b��<���<G��<]��<G��<���<b��<@��<c��<���<�	�<7�<�%�<`0�<v7�<`   `   	?�<5=�<�5�<i*�<_�<��<��<\��<:��<e��<��<x��<S��<x��<��<e��<:��<\��<��<��<_�<i*�<�5�<5=�<`   `   �@�<�>�<47�<�+�<q�<�<T��<���<:��<}��<���<Q��<��<Q��<���<}��<:��<���<T��<�<q�<�+�<47�<�>�<`   `   >?�<+<�<l4�<�(�<�<��<t��<��<���<���<���< ��<r��< ��<���<���<���<��<t��<��<�<�(�<l4�<+<�<`   `   
:�<+7�</�<�"�<I�<p�<��<t��<h��<e��<=��<ަ�<��<ަ�<=��<e��<h��<t��<��<p�<I�<�"�</�<+7�<`   `   y0�<t.�<�&�<��<e�<W��<���<���<��<���<d��<���<W��<���<d��<���<��<���<���<W��<e�<��<�&�<t.�<`   `   I%�<W#�<��<�<H�<���<���<��<���<!��<���<���<���<���<���<!��<���<��<���<���<H�<�<��<W#�<`   `   i�<�<��<��<��<��<!��< ��<:��< ��<���<���<���<���<���< ��<:��< ��<!��<��<��<��<��<�<`   `   ��<=	�<i�<���<?��<1��<X��<ظ�<���<F��<���<��<���<��<���<F��<���<ظ�<X��<1��<?��<���<i�<=	�<`   `   l��<_��<0��<���<���<:��<R��<z��<��<���<5��<*��<.��<*��<5��<���<��<z��<R��<:��<���<���<0��<_��<`   `   ���< ��<���<|��<���<���<��<���<w��<���<��<���<��<���<��<���<w��<���<��<���<���<|��<���< ��<`   `   ���<���<F��<H��<o��<&��<ӳ�<��<h��<3��<^��<���<D��<���<^��<3��<h��<��<ӳ�<&��<o��<H��<F��<���<`   `   ���<���<?��<���<���<���<���<���<��<z��<��<��<ǉ�<��<��<z��<��<���<���<���<���<���<?��<���<`   `   ���<+��<G��<y��<���<��<��<���<���</��<v��<v��<D��<v��<v��</��<���<���<��<��<���<y��<G��<+��<`   `   ���<���<6��<���<��<e��<���<ʫ�<���<.��<���<���<|��<���<���<.��<���<ʫ�<���<e��<��<���<6��<���<`   `   .��<���<5��<i��<���<"��< ��<a��<���<���<��<���<���<���<��<���<���<a��< ��<"��<���<i��<5��<���<`   `   )��<���<U��<(��<H��<#��<U��<Ϻ�<0��<~��<>��<5��<���<5��<>��<~��<0��<Ϻ�<U��<#��<H��<(��<U��<���<`   `   ���<��<'��<��<W��<���<��<_��<p��<T��<@��<U��<t��<U��<@��<T��<p��<_��<��<���<W��<��<'��<��<`   `   Խ�<���<9��<5��<���<���<>��<��<e��<S��<���<���<@��<���<���<S��<e��<��<>��<���<���<5��<9��<���<`   `   ���<���<���<���<���<���<��<.��<���<L��<���<��<���<��<���<L��<���<.��<��<���<���<���<���<���<`   `   y��</��<Q��<T��<��<���<���<���<"��<t��<Q��<��<�<��<Q��<t��<"��<���<���<���<��<T��<Q��</��<`   `   ���<���<���<���<���<N��<6��<\��<e��<�<J�<u�<�<u�<J�<�<e��<\��<6��<N��<���<���<���<���<`   `   p��<���<���<9��<y��<���<_��<|��<�	�<y�<��<�!�<V#�<�!�<��<y�<�	�<|��<_��<���<y��<9��<���<���<`   `   O��<��<���<J��<���<���<0��<�<�<��<7(�<U.�<�/�<U.�<7(�<��<�<�<0��<���<���<J��<���<��<`   `   ]��<G��<���<b��<@��<c��<���<�	�<7�<�%�<`0�<v7�<�8�<v7�<`0�<�%�<7�<�	�<���<c��<@��<b��<���<G��<`   `   S��<x��<��<e��<:��<\��<��<��<_�<i*�<�5�<5=�<	?�<5=�<�5�<i*�<_�<��<��<\��<:��<e��<��<x��<`   `   ��<Q��<���<}��<:��<���<T��<�<q�<�+�<47�<�>�<�@�<�>�<47�<�+�<q�<�<T��<���<:��<}��<���<Q��<`   `   r��< ��<���<���<���<��<t��<��<�<�(�<l4�<+<�<>?�<+<�<l4�<�(�<�<��<t��<��<���<���<���< ��<`   `   ��<ަ�<=��<e��<h��<t��<��<p�<I�<�"�</�<+7�<
:�<+7�</�<�"�<I�<p�<��<t��<h��<e��<=��<ަ�<`   `   W��<���<d��<���<��<���<���<W��<f�<��<�&�<t.�<y0�<t.�<�&�<��<f�<W��<���<���<��<���<d��<���<`   `   ���<���<���<!��<���<��<���<���<H�< �<��<W#�<I%�<W#�<��< �<H�<���<���<��<���<!��<���<���<`   `   ���<���<���< ��<:��< ��<!��<��<��<��<��<�<j�<�<��<��<��<��<!��< ��<:��< ��<���<���<`   `   ���<��<���<F��<���<ظ�<X��<1��<?��<���<i�<=	�<��<=	�<i�<���<?��<1��<X��<ظ�<���<F��<���<��<`   `   .��<*��<5��<���<��<z��<R��<:��<���<���<0��<_��<l��<_��<0��<���<���<:��<R��<z��<��<���<5��<*��<`   `   �j�<zm�<]t�<��<i��<���<���<y��<P��<���<K��<���<=��<���<K��<���<P��<y��<���<���<i��<��<]t�<zm�<`   `   �l�<o�<u�<�~�<���<���<6��<o��<(��<f��<���<4��<0��<4��<���<f��<(��<o��<6��<���<���<�~�<u�<o�<`   `   s�<�t�<ny�<ȁ�<���<1��<��<���<���<���<B��<��<���<��<B��<���<���<���<��<1��<���<ȁ�<ny�<�t�<`   `   �|�<~�<��<���<h��<0��<��<а�<%��<���<h��<��<��<��<h��<���<%��<а�<��<0��<h��<���<��<~�<`   `   ��<��<Ɏ�<A��<q��<���<H��<Ư�<_��<���<���<��<���<��<���<���<_��<Ư�<H��<���<q��<A��<Ɏ�<��<`   `   <��<z��<���<k��<��<x��<ӭ�<K��<۶�<���<��<��<L��<��<��<���<۶�<K��<ӭ�<x��<��<k��<���<z��<`   `   K��<��<H��<I��<��<��<B��<���<���<3��<x��<'��<���<'��<x��<3��<���<���<B��<��<��<I��<H��<��<`   `   ���<`��<���<X��< ��<-��<*��<��<A��<+��<��<��<d��<��<��<+��<A��<��<*��<-��< ��<X��<���<`��<`   `   ���<6��<&��<���< ��<��<n��<���<7��<���<\��<4��<���<4��<\��<���<7��<���<n��<��< ��<���<&��<6��<`   `   n��<b��<��<p��<���<:��<=��<���<���<a��<���<w��<���<w��<���<a��<���<���<=��<:��<���<p��<��<b��<`   `   ��<.�<��<0�<���<��<7��<���<���<;��<���<���<���<���<���<;��<���<���<7��<��<���<0�<��<.�<`   `   �-�<g+�<�%�<k�< �<��<��<z��<���</��<���<|��<��<|��<���</��<���<z��<��<��< �<k�<�%�<g+�<`   `   �B�<�?�<�8�<�-�<m�<�<>��<���<���<���<n��<��<���<��<n��<���<���<���<>��<�<m�<�-�<�8�<�?�<`   `   {S�<�P�<�H�<<�<�+�<��<��<���<���<���<}��<<��<���<<��<}��<���<���<���<��<��<�+�<<�<�H�<�P�<`   `   �_�<�\�<XT�<F�<4�<>�<		�<���<���<p��<`��<���<��<���<`��<p��<���<���<		�<>�<4�<F�<XT�<�\�<`   `   Gg�<�c�<�Z�<:L�<�8�<A"�<Y
�<���<���<	��<���<���<���<���<���<	��<���<���<Y
�<A"�<�8�<:L�<�Z�<�c�<`   `   9j�<Nf�<�\�<
M�<N8�<'!�<��<��<���<��<C��<��<���<��<C��<��<���<��<��<'!�<N8�<
M�<�\�<Nf�<`   `   �f�<�c�<�Y�<�I�<J4�<�<�<q��<���<���<���<L��<��<L��<���<���<���<q��<�<�<J4�<�I�<�Y�<�c�<`   `   f_�<W\�<\R�<B�<�,�<��<���<���<���<&��<P��<���<"��<���<P��<&��<���<���<���<��<�,�<B�<\R�<W\�<`   `   �T�<2Q�<�F�<d6�<_!�<~�<���<��<���<I��<Θ�<`��< ��<`��<Θ�<I��<���<��<���<~�<_!�<d6�<�F�<2Q�<`   `   �E�< B�<�7�<(�<e�<���<D��<��<���<ŝ�<���<���<��<���<���<ŝ�<���<��<D��<���<e�<(�<�7�< B�<`   `   &4�<�0�<�'�<n�<\�<���<3��</��<��<��<$��<�{�<�x�<�{�<$��<��<��</��<3��<���<\�<n�<�'�<�0�<`   `   �!�<Z�<��<X�<���<i��<_��<���<��<ъ�<}�<{t�<�q�<{t�<}�<ъ�<��<���<_��<i��<���<X�<��<Z�<`   `   ��<��<��<t��<5��<���<���<H��<X��<���<5w�<�o�<�l�<�o�<5w�<���<X��<H��<���<���<5��<t��<��<��<`   `   <��<���<K��<���<P��<y��<���<���<i��<��<]t�<zm�<�j�<zm�<]t�<��<i��<���<���<y��<P��<���<K��<���<`   `   0��<4��<���<f��<(��<o��<6��<���<���<�~�<u�<o�<�l�<o�<u�<�~�<���<���<6��<o��<(��<f��<���<4��<`   `   ���<��<B��<���<���<���<��<1��<���<ȁ�<my�<�t�<s�<�t�<my�<ȁ�<���<1��<��<���<���<���<B��<��<`   `   ��<��<h��<���<%��<а�<��<0��<h��<���<��<~�<�|�<~�<��<���<h��<0��<��<а�<%��<���<h��<��<`   `   ���<��<���<���<_��<Ư�<H��<���<q��<A��<Ɏ�<��<��<��<Ɏ�<A��<q��<���<H��<Ư�<_��<���<���<��<`   `   L��<��<��<���<۶�<K��<ӭ�<x��<��<k��<���<z��<;��<z��<���<k��<��<x��<ӭ�<K��<۶�<���<��<��<`   `   ���<'��<x��<3��<���<���<B��<��<��<I��<G��<��<K��<��<G��<I��<��<��<B��<���<���<3��<x��<'��<`   `   d��<��<��<+��<A��<��<*��<-��< ��<X��<���<`��<���<`��<���<X��< ��<-��<*��<��<A��<+��<��<��<`   `   ���<4��<\��<���<7��<���<n��<��< ��<���<&��<6��<���<6��<&��<���< ��<��<n��<���<7��<���<\��<4��<`   `   ���<w��<���<a��<���<���<=��<:��<���<p��<��<b��<n��<b��<��<p��<���<:��<=��<���<���<a��<���<w��<`   `   ���<���<���<;��<���<���<7��<��<���<0�<��<.�<��<.�<��<0�<���<��<7��<���<���<;��<���<���<`   `   ��<|��<���</��<���<z��<��<��< �<k�<�%�<g+�<�-�<g+�<�%�<k�< �<��<��<z��<���</��<���<|��<`   `   ���<��<n��<���<���<���<>��<�<m�<�-�<�8�<�?�<�B�<�?�<�8�<�-�<m�<�<>��<���<���<���<n��<��<`   `   ���<<��<~��<���<���<���<��<��<�+�<<�<�H�<�P�<{S�<�P�<�H�<<�<�+�<��<��<���<���<���<}��<<��<`   `   ��<���<`��<p��<���<���<		�<>�<4�<F�<XT�<�\�<�_�<�\�<XT�<F�<4�<>�<		�<���<���<p��<`��<���<`   `   ���<���<���<	��<���<���<Y
�<A"�<�8�<:L�<�Z�<�c�<Gg�<�c�<�Z�<:L�<�8�<A"�<Y
�<���<���<	��<���<���<`   `   ���<��<C��<��<���<��<��<'!�<N8�<
M�<�\�<Nf�<9j�<Nf�<�\�<
M�<N8�<'!�<��<��<���<��<C��<��<`   `   ��<L��<���<���<���<q��<�<�<J4�<�I�<�Y�<�c�<�f�<�c�<�Y�<�I�<J4�<�<�<q��<���<���<���<L��<`   `   "��<���<P��<&��<���<���<���<��<�,�<B�<\R�<W\�<f_�<W\�<\R�<B�<�,�<��<���<���<���<&��<P��<���<`   `    ��<`��<Θ�<I��<���<��<���<~�<_!�<e6�<�F�<2Q�<�T�<2Q�<�F�<e6�<_!�<~�<���<��<���<I��<Θ�<`��<`   `   ��<���<���<ŝ�<���<��<D��<���<f�<(�<�7�< B�<�E�< B�<�7�<(�<f�<���<D��<��<���<ŝ�<���<���<`   `   �x�<�{�<$��<��<��</��<3��<���<\�<o�<�'�<�0�<&4�<�0�<�'�<o�<\�<���<3��</��<��<��<$��<�{�<`   `   �q�<{t�<}�<ъ�<��<���<_��<i��<���<X�<��<Z�<�!�<Z�<��<X�<���<i��<_��<���<��<ъ�<}�<{t�<`   `   �l�<�o�<5w�<���<X��<H��<���<���<5��<u��<��<��<��<��<��<u��<5��<���<���<H��<X��<���<5w�<�o�<`   `   &H�<�K�<�T�<d�<\x�<���<ި�<;��<E��<g��<���<f�<��<f�<���<g��<E��<;��<ި�<���<\x�<d�<�T�<�K�<`   `   �J�<�M�<DV�<�b�<�t�<���<���<y��<j��<R��<���<T��<���<T��<���<R��<j��<y��<���<���<�t�<�b�<DV�<�M�<`   `   �R�<U�<5\�<�f�<wu�<!��<y��<m��<��<���<k��<��<���<��<k��<���<��<m��<y��<!��<wu�<�f�<5\�<U�<`   `   &`�<�a�<�g�<p�<�{�<���</��<��<���<ڿ�<��<6��<���<6��<��<ڿ�<���<��</��<���<�{�<p�<�g�<�a�<`   `   Hs�<xt�<�x�<�~�<|��<��<���<S��<%��<��<���<��<}��<��<���<��<%��<S��<���<��<|��<�~�<�x�<xt�<`   `   :��<Ӌ�<���<ޑ�<,��<
��<��<���<ޮ�<ֳ�<���<d��<E��<d��<���<ֳ�<ޮ�<���<��<
��<,��<ޑ�<���<Ӌ�<`   `   ���<���<���<s��<s��<+��<6��<���<w��<���<��<D��<���<D��<��<���<w��<���<6��<+��<s��<s��<���<���<`   `   a��<���<���<���<���<��<��<���<c��<���<���<C��<���<C��<���<���<c��<���<��<��<���<���<���<���<`   `   ���<���<c��<���<��<���<���<���<^��<��<���<Y��<:��<Y��<���<��<^��<���<���<���<��<���<c��<���<`   `   ��<�
�<��<���<��<���< ��<���<���<���<��<}��<[��<}��<��<���<���<���< ��<���<��<���<��<�
�<`   `   O.�<',�<�%�<a�<��<9��<���<Q��<���<d��<»�<��<��<��<»�<d��<���<Q��<���<9��<��<a�<�%�<',�<`   `   dN�<�K�<�C�<k6�<`&�<|�<���<���<S��<b��<_��<B��<δ�<B��<_��<b��<S��<���<���<|�<`&�<k6�<�C�<�K�<`   `   lj�</g�<�]�<�N�<T;�<�$�<9�<���< ��<���<~��<��<���<��<~��<���< ��<���<9�<�$�<T;�<�N�<�]�</g�<`   `   ā�<�}�<s�<�a�<�K�<'2�<E�<A��<��<���<w��<���<���<���<w��<���<��<A��<E�<'2�<�K�<�a�<s�<�}�<`   `   ���<���<��<p�<aW�<;�<�<4��<���<���<��<0��<���<0��<��<���<���<4��<�<;�<aW�<p�<��<���<`   `   ܝ�<ژ�<���<�w�<I]�<�>�<l�<���<:��<��<˴�<Ȩ�< ��<Ȩ�<˴�<��<:��<���<l�<�>�<I]�<�w�<���<ژ�<`   `   z��<g��<���<�x�<Y]�<P=�<�<���<��<��<%��<Z��<(��<Z��<$��<��<��<���<�<P=�<Y]�<�x�<���<g��<`   `   ���<��<���<"t�<X�<�6�<��<���<V��<���<��<���<a��<���<��<���<V��<���<��<�6�<X�<"t�<���<��<`   `   ��<8��<��<�i�<�L�<�+�<5�<���<���<<��<���<���<��<���<���<<��<���<���<5�<�+�<�L�<�i�<��<8��<`   `   t��<Z~�<]p�<wZ�<�=�<��<���<l��<~��<7��<^��<Jy�<�t�<Jy�<^��<7��<~��<l��<���<��<�=�<wZ�<]p�<Z~�<`   `   Bo�<Aj�<�\�<�G�<3+�<d�<���<���<O��<���<�x�<�k�<�f�<�k�<�x�<���<O��<���<���<d�<3+�<�G�<�\�<Aj�<`   `   �W�<S�<F�<.1�<��<���<���<���<\��<�~�<Sk�<_�<8[�<_�<Sk�<�~�<\��<���<���<���<��<.1�<F�<S�<`   `   >�<:�<�-�<7�<{�<���<���<��<ފ�<�r�<p`�<"U�<�Q�<"U�<p`�<�r�<ފ�<��<���<���<{�<7�<�-�<:�<`   `   �$�<� �<]�<�<���<���<��<���<��<�i�<�X�<\N�<�J�<\N�<�X�<�i�<��<���<��<���<���<�<]�<� �<`   `   ��<e�<���<g��<E��<:��<ި�<���<\x�<d�<�T�<�K�<&H�<�K�<�T�<d�<\x�<���<ި�<:��<E��<g��<���<e�<`   `   ���<T��<���<R��<j��<y��<���<���<�t�<�b�<DV�<�M�<�J�<�M�<DV�<�b�<�t�<���<���<y��<j��<R��<���<T��<`   `   ���<��<k��<���<��<m��<y��<!��<wu�<�f�<5\�<U�<�R�<U�<5\�<�f�<wu�<!��<y��<m��<��<���<k��<��<`   `   ���<6��<��<ڿ�<���<��</��<���<�{�<p�<�g�<�a�<&`�<�a�<�g�<p�<�{�<���</��<��<���<ڿ�<��<6��<`   `   }��<��<���<��<%��<S��<���<��<|��<�~�<�x�<xt�<Hs�<xt�<�x�<�~�<|��<��<���<S��<%��<��<���<��<`   `   E��<c��<���<ֳ�<ޮ�<���<��<	��<,��<ޑ�<���<Ӌ�<:��<Ӌ�<���<ޑ�<,��<	��<��<���<ޮ�<ֳ�<���<c��<`   `   ���<D��<��<���<w��<���<5��<+��<r��<s��<���<���<���<���<���<s��<r��<+��<5��<���<w��<���<��<D��<`   `   ���<C��<���<���<c��<���<��<��<���<���<���<���<a��<���<���<���<���<��<��<���<c��<���<���<C��<`   `   :��<Y��<���<��<^��<���<���<���<��<���<c��<���<���<���<c��<���<��<���<���<���<^��<��<���<Y��<`   `   [��<}��<��<���<���<���< ��<���<��<���<��<�
�<��<�
�<��<���<��<���< ��<���<���<���<��<}��<`   `   ��<��<»�<d��<���<Q��<���<9��<��<a�<�%�<',�<O.�<',�<�%�<a�<��<9��<���<Q��<���<d��<»�<��<`   `   δ�<B��<_��<b��<S��<���<���<|�<`&�<k6�<�C�<�K�<dN�<�K�<�C�<k6�<`&�<|�<���<���<S��<b��<_��<B��<`   `   ���<��<~��<���< ��<���<9�<�$�<T;�<�N�<�]�</g�<lj�</g�<�]�<�N�<T;�<�$�<9�<���< ��<���<~��<��<`   `   ���<���<w��<���<��<A��<E�<'2�<�K�<�a�<s�<�}�<ā�<�}�<s�<�a�<�K�<'2�<E�<A��<��<���<w��<���<`   `   ���<0��<��<���<���<4��<�<;�<aW�<p�<��<���<���<���<��<p�<aW�<;�<�<4��<���<���<��<0��<`   `    ��<Ȩ�<˴�<��<:��<���<l�<�>�<I]�<�w�<���<ژ�<ܝ�<ژ�<���<�w�<I]�<�>�<l�<���<:��<��<˴�<Ȩ�<`   `   (��<Z��<%��<��<��<���<�<Q=�<Y]�<�x�<���<g��<z��<g��<���<�x�<Y]�<Q=�<�<���<��<��<%��<Z��<`   `   a��<���<��<���<V��<���<��<�6�<X�<"t�<���<��<���<��<���<"t�<X�<�6�<��<���<V��<���<��<���<`   `   ��<���<���<<��<���<���<5�<�+�<�L�<�i�<��<8��<��<8��<��<�i�<�L�<�+�<5�<���<���<<��<���<���<`   `   �t�<Ky�<^��<7��<~��<l��<���<��<�=�<wZ�<]p�<Z~�<u��<Z~�<]p�<wZ�<�=�<��<���<l��<~��<7��<^��<Jy�<`   `   �f�<�k�<�x�<���<O��<���<���<e�<3+�<�G�<�\�<Bj�<Bo�<Bj�<�\�<�G�<3+�<e�<���<���<O��<���<�x�<�k�<`   `   8[�<_�<Sk�<�~�<\��<���<���<���<��<.1�<F�<S�<�W�<S�<F�<.1�<��<���<���<���<\��<�~�<Sk�<_�<`   `   �Q�<"U�<p`�<�r�<ފ�<��<���<���<{�<7�<�-�<:�<>�<:�<�-�<7�<{�<���<���<��<ފ�<�r�<p`�<"U�<`   `   �J�<\N�<�X�<�i�<��<���<��<���<���<�<]�<� �<�$�<� �<]�<�<���<���<��<���<��<�i�<�X�<\N�<`   `   ~�<*�<�)�<>�<VX�<:w�<��<��<	��<m��<[�<��<�<��<[�<m��<��<��<��<:w�<UX�<>�<�)�<*�<`   `   ��<��<+�<�<�<�S�<�n�<��<=��<���<4��<��<���<� �<���<��<4��<���<=��<��<�n�<�S�<�<�<+�<��<`   `   ('�<�)�<�3�<�A�<�T�<�k�<j��<D��<]��<Z��<���<���<:��<���<���<Z��<]��<D��<j��<�k�<�T�<�A�<�3�<�)�<`   `   �9�<m;�<�B�<�M�<N]�<Co�<҂�<m��<���<{��<|��<��<���<��<|��<{��<���<m��<҂�<Co�<N]�<�M�<�B�<m;�<`   `   �R�<�S�<�X�<#a�<;l�<�x�<��<F��<���<��<���<���<��<���<���<��<���<F��<��<�x�<;l�<#a�<�X�<�S�<`   `   =r�<-s�<v�<�z�<:��<���<F��<���<ӡ�<j��<���<z��<T��<z��<���<j��<ӡ�<���<F��<���<:��<�z�<v�<-s�<`   `   ���<��<1��<��<��<��<P��<��<��<���<Ԫ�<2��<4��<2��<Ԫ�<���<��<��<P��<��<��<��<1��<��<`   `   O��<���<���<���<���<���<̳�< ��<8��<ū�<���<s��<��<s��<���<ū�<8��< ��<̳�<���<���<���<���<���<`   `   ���<���<m��<���<���<��<\��<��<���<J��<���<`��<��<`��<���<J��<���<��<\��<��<���<���<m��<���<`   `   k �</�<��<��<G �<���<��<>��<���<��<���<6��<��<6��<���<��<���<>��<��<���<G �<��<��</�<`   `   |N�<�K�<�B�<�4�<#�<�<���<��<��<F��<���<��<x��<��<���<F��<��<��<���<�<#�<�4�<�B�<�K�<`   `   �y�<v�<Ck�<�Y�<�C�<#*�<��<'��<���<l��<L��<խ�<���<խ�<L��<l��<���<'��<��<#*�<�C�<�Y�<Ck�<v�<`   `   Q��<��<��<xz�<`�<A�<� �<k�</��<~��<ո�<g��<f��<g��<ո�<~��</��<k�<� �<A�<`�<xz�<��<��<`   `   ���<ں�<���<���<�v�<iS�<�.�<�
�<0��<���<ܷ�<Z��<T��<Z��<ܷ�<���<0��<�
�<�.�<iS�<�v�<���<���<ں�<`   `   ��<���<k��<5��<G��<�_�<(7�<��<���<���<���<ӣ�<���<ӣ�<���<���<���<��<(7�<�_�<G��<5��<k��<���<`   `   "��<���<R��<
��<*��<�d�<�8�<C�<���<��<��<
��<۔�<
��<��<��<���<C�<�8�<�d�<*��<
��<R��<���<`   `   R��<z��<���<L��<a��<�b�<c4�<��<.��<���<M��<��<�<��<M��<���<.��<��<c4�<�b�<a��<L��<���<z��<`   `   ���<���<���<���<ۆ�<�Y�<f*�<���<X��<���<o��<~�< x�<~�<o��<���<X��<���<f*�<�Y�<ۆ�<���<���<���<`   `   ���</��<���<3��<�w�<�J�<��<���<+��<	��<�}�<il�<of�<il�<�}�<	��<+��<���<��<�J�<�w�<3��<���</��<`   `   ���<���<���<n��<&c�<o6�<��<g��<N��<*��<7k�<�Y�<�S�<�Y�<7k�<*��<N��<g��<��<o6�<&c�<n��<���<���<`   `   ��<���<t��<,p�<9J�<��<���<���<n��<t�<�X�<�G�<�A�<�G�<�X�<t�<n��<���<���<��<9J�<,p�<t��<���<`   `   8��<a��<{n�<KR�<t.�<e�<!��<Ƭ�<���<�a�<�G�<�7�<Q2�<�7�<�G�<�a�<���<Ƭ�<!��<e�<t.�<KR�<{n�<a��<`   `   �c�<n^�<�M�<43�<��<)��<���<'��<�q�<�Q�<�9�<�)�<X$�<�)�<�9�<�Q�<�q�<'��<���<)��<��<43�<�M�<n^�<`   `   �@�<�;�<�,�<Y�<���<���<��<���<�b�<�E�<//�<� �<��<� �<//�<�E�<�b�<���<��<���<���<Y�<�,�<�;�<`   `   �<��<[�<m��<��<��<��<:w�<UX�<>�<�)�<*�<}�<*�<�)�<>�<UX�<:w�<��<��<��<m��<[�<��<`   `   � �<���<��<3��<���<=��< ��<�n�<�S�<�<�<+�<��<��<��<+�<�<�<�S�<�n�< ��<=��<���<3��<��<���<`   `   :��<���<���<Z��<]��<D��<j��<�k�<�T�<�A�<�3�<�)�<('�<�)�<�3�<�A�<�T�<�k�<j��<D��<]��<Z��<���<���<`   `   ���<��<|��<z��<���<m��<т�<Bo�<N]�<�M�<�B�<m;�<�9�<m;�<�B�<�M�<N]�<Bo�<т�<m��<���<z��<|��<��<`   `   ��<���<���<��<���<F��<��<�x�<;l�<#a�<�X�<�S�<�R�<�S�<�X�<#a�<;l�<�x�<��<F��<���<��<���<���<`   `   T��<z��<���<j��<ӡ�<���<F��<���<:��<�z�<v�<-s�<=r�<-s�<v�<�z�<:��<���<F��<���<ӡ�<j��<���<z��<`   `   4��<2��<Ԫ�<���<��<��<P��<��<��<��<1��<��<���<��<1��<��<��<��<P��<��<��<���<Ԫ�<2��<`   `   ��<s��<���<ū�<8��< ��<̳�<���<���<���<���<���<O��<���<���<���<���<���<̳�< ��<8��<ū�<���<s��<`   `   ��<_��<���<J��<���<��<\��<��<���<���<m��<���<���<���<m��<���<���<��<\��<��<���<J��<���<_��<`   `   ��<6��<���<��<���<>��<��<���<G �<��<��</�<k �</�<��<��<G �<���<��<>��<���<��<���<6��<`   `   x��<��<���<F��<��<��<���<�<#�<�4�<�B�<�K�<|N�<�K�<�B�<�4�<#�<�<���<��<��<F��<���<��<`   `   ���<խ�<L��<l��<���<'��<��<#*�<�C�<�Y�<Ck�<v�<�y�<v�<Ck�<�Y�<�C�<#*�<��<'��<���<l��<L��<խ�<`   `   f��<g��<ո�<~��</��<k�<� �<A�<`�<xz�<��<��<Q��<��<��<xz�<`�<A�<� �<k�</��<~��<ո�<g��<`   `   T��<Z��<ܷ�<���<0��<�
�<�.�<iS�<�v�<���<���<ں�<���<ں�<���<���<�v�<iS�<�.�<�
�<0��<���<ܷ�<Z��<`   `   ���<ӣ�<���<���<���<��<(7�<�_�<G��<5��<k��<���<��<���<k��<5��<G��<�_�<(7�<��<���<���<���<ӣ�<`   `   ۔�<
��<��<��<���<C�<�8�<�d�<+��<
��<R��<���<"��<���<R��<
��<+��<�d�<�8�<C�<���<��<��<
��<`   `   �<��<M��<���</��<��<c4�<�b�<a��<L��<���<z��<R��<z��<���<L��<a��<�b�<c4�<��<.��<���<M��<��<`   `    x�<~�<o��<���<X��<���<f*�<�Y�<ۆ�<���<���<���<���<���<���<���<ۆ�<�Y�<f*�<���<X��<���<o��<~�<`   `   of�<il�<�}�<	��<+��<���<��<�J�<�w�<3��<���</��<���</��<���<3��<�w�<�J�<��<���<+��<	��<�}�<il�<`   `   �S�<�Y�<7k�<*��<N��<h��<��<p6�<'c�<n��<���<���<���<���<���<n��<'c�<p6�<��<g��<N��<*��<7k�<�Y�<`   `   �A�<�G�<�X�<t�<n��<���<���<��<9J�<,p�<t��<���<��<���<t��<,p�<9J�<��<���<���<n��<t�<�X�<�G�<`   `   Q2�<�7�<�G�<�a�<���<Ƭ�<!��<e�<t.�<KR�<{n�<a��<8��<a��<{n�<KR�<t.�<e�<!��<Ƭ�<���<�a�<�G�<�7�<`   `   X$�<�)�<�9�<�Q�<�q�<'��<���<)��<��<43�<�M�<n^�<�c�<n^�<�M�<43�<��<)��<���<'��<�q�<�Q�<�9�<�)�<`   `   ��<� �<//�<�E�<�b�<���<��<���<���<Y�<�,�<�;�<�@�<�;�<�,�<Y�<���<���<��<���<�b�<�E�<//�<� �<`   `   ���<K��<��<�	�< -�<7W�<��<��<��<��<
 �<52�<�8�<52�<
 �<��<��<��<��<7W�< -�<�	�<��<K��<`   `   T��<���<b��<��<�&�<CK�<r�<ۙ�<���<���<���<�	�<��<�	�<���<���<���<ۙ�<r�<CK�<�&�<��<b��<���<`   `   ?��<��<@��<��<u(�<	G�<�g�<��<ڨ�<[��<���<.��<`��<.��<���<[��<ڨ�<��<�g�<	G�<u(�<��<@��<��<`   `   n�<��<��<�<R3�<AK�<he�<���<ƙ�< ��<J��<0��<���<0��<J��< ��<ƙ�<���<he�<AK�<R3�<�<��<��<`   `   �$�<'�<�-�< 9�<G�<cX�<$k�<�~�<\��<נ�<��< ��<���< ��<��<נ�<\��<�~�<$k�<cX�<G�< 9�<�-�<'�<`   `   �O�<8Q�<U�<�[�<�c�<�m�<|y�<��<r��<X��<y��<{��<z��<{��<y��<X��<r��<��<|y�<�m�<�c�<�[�<U�<8Q�<`   `   &��<���<Ƀ�<J��<1��<��<���<��<��<��<���<���<c��<���<���<��<��<��<���<��<1��<J��<Ƀ�<���<`   `   ۻ�<���<0��<���<-��<B��<7��<���<���<��<��<��<Ú�<��<��<��<���<���<7��<B��<-��<���<0��<���<`   `   ���<6��<���<���<���<���<��<й�<\��<5��<?��<,��<���<,��<?��<5��<\��<й�<��<���<���<���<���<6��<`   `   j9�<�6�<�-�<��<6�<���<���<���<���<¯�<<��<,��<���<,��<<��<¯�<���<���<���<���<6�<��<�-�<�6�<`   `   �x�<Pt�<�h�<V�<�=�<)"�</�<`��<���<|��<���<���<��<���<���<|��<���<`��</�<)"�<�=�<V�<�h�<Pt�<`   `   ���<��<��<܇�<Ii�<�F�<\"�< ��<t��<���<\��<$��<m��<$��<\��<���<t��< ��<\"�<�F�<Ii�<܇�<��<��<`   `   ��<���<s��<���<G��<�f�<8;�<q�<��<k��<ͯ�<��<���<��<ͯ�<k��<��<q�<8;�<�f�<G��<���<s��<���<`   `   �<�<���<���<f��<X�<CM�<)�<���<���<��<2��<v��<2��<��<���<���<)�<CM�<X�<f��<���<���<�<`   `   �2�<H+�<��<���<���<1��<X�<�!�<U��<=��<o��<���<��<���<o��<=��<U��<�!�<X�<1��<���<���<��<H+�<`   `   #G�<�>�<�%�< �<���<Z��</[�<H �<���<#��<=��<܅�<#~�<܅�<=��<#��<���<H �</[�<Z��<���< �<�%�<�>�<`   `   �M�<�D�<�*�<��<���<ȓ�<RU�<�<���<���<���<Pt�<(l�<Pt�<���<���<���<�<RU�<ȓ�<���<��<�*�<�D�<`   `   �F�<a=�<#�<���<e��<k��<�F�<4�<B��<���<3v�<_�<�V�<_�<3v�<���<B��<4�<�F�<k��<e��<���<#�<a=�<`   `   3�<)*�<�<���<Ȱ�<s�<�1�<���<ܶ�<��<�_�<�G�<�?�<�G�<�_�<��<ܶ�<���<�1�<s�<Ȱ�<���<�<)*�<`   `   ��<��<���<���<Ĕ�<�W�<*�<���<g��<l�<�F�<'/�<6'�<'/�<�F�<l�<g��<���<*�<�W�<Ĕ�<���<���<��<`   `   ��<V��<���<���<]r�<7�<{��<���<��<;R�<�-�<��<�<��<�-�<;R�<��<���<{��<7�<]r�<���<���<V��<`   `   ��<���<���<�}�<�L�<>�<���<���<.g�<�9�<��<� �<g��<� �<��<�9�<.g�<���<���<>�<�L�<�}�<���<���<`   `   ��<��<w�<�S�<n%�<���<8��<���<'O�<$�<!�<���<���<���<!�<$�<'O�<���<8��<���<n%�<�S�<w�<��<`   `   Df�<�^�<3J�<�)�<I��<@��<��<�i�<<;�<R�<���<-��<���<-��<���<R�<<;�<�i�<��<@��<I��<�)�<3J�<�^�<`   `   �8�<42�<
 �<��<��<��<��<6W�< -�<�	�<��<K��<���<K��<��<�	�< -�<6W�<��<��<��<��<
 �<42�<`   `   ��<�	�<���<���<���<ۙ�<r�<BK�<�&�<��<b��<���<S��<���<b��<��<�&�<BK�<r�<ۙ�<���<���<���<�	�<`   `   `��<.��<���<[��<ڨ�<��<�g�<	G�<u(�<��<@��<��<?��<��<@��<��<u(�<	G�<�g�<��<ڨ�<[��<���<.��<`   `   ���<0��<J��< ��<ƙ�<���<he�<AK�<R3�<�<��<��<n�<��<��<�<R3�<AK�<he�<���<ƙ�< ��<J��<0��<`   `   ���<���<��<נ�<\��<�~�<#k�<cX�<~G�< 9�<�-�<'�<�$�<'�<�-�< 9�<~G�<cX�<#k�<�~�<\��<נ�<��<���<`   `   z��<{��<y��<X��<q��<��<{y�<�m�<�c�<�[�<U�<7Q�<�O�<7Q�<U�<�[�<�c�<�m�<{y�<��<q��<X��<y��<{��<`   `   c��<���<���<��<��<��<���<��<1��<J��<Ƀ�<���<&��<���<Ƀ�<J��<1��<��<���<��<��<��<���<���<`   `   Ú�<��<��<��<���<���<7��<B��<-��<���<0��<���<ۻ�<���<0��<���<-��<B��<7��<���<���<��<��<��<`   `   ���<+��<?��<5��<\��<й�<��<���<���<���<���<6��<���<6��<���<���<���<���<��<й�<\��<5��<?��<+��<`   `   ���<,��<;��<¯�<���<���<���<���<6�<��<�-�<�6�<j9�<�6�<�-�<��<6�<���<���<���<���<¯�<;��<,��<`   `   ��<���<���<|��<���<`��</�<)"�<�=�<V�<�h�<Pt�<�x�<Pt�<�h�<V�<�=�<)"�</�<`��<���<|��<���<���<`   `   m��<$��<\��<���<t��< ��<\"�<�F�<Ii�<܇�<��<��<���<��<��<܇�<Ii�<�F�<\"�< ��<t��<���<\��<$��<`   `   ���<��<ͯ�<k��<��<q�<8;�<�f�<G��<���<s��<���<��<���<s��<���<G��<�f�<8;�<q�<��<k��<ͯ�<��<`   `   v��<2��<��<���<���<)�<CM�<X�<f��<���<���<�<�<�<���<���<f��<X�<CM�<)�<���<���<��<2��<`   `   ��<���<o��<=��<U��<�!�<X�<1��<���<���<��<H+�<�2�<H+�<��<���<���<1��<X�<�!�<U��<=��<o��<���<`   `   #~�<܅�<=��<#��<���<H �</[�<Z��<���< �<�%�<�>�<#G�<�>�<�%�< �<���<Z��</[�<H �<���<#��<=��<܅�<`   `   (l�<Qt�<���<���<���<�<RU�<ȓ�<���<��<�*�<�D�<�M�<�D�<�*�<��<���<ȓ�<RU�<�<���<���<���<Qt�<`   `   �V�<_�<3v�<���<B��<4�<�F�<k��<e��<���<#�<a=�<�F�<a=�<#�<���<e��<k��<�F�<4�<B��<���<3v�<_�<`   `   �?�<�G�<�_�<��<ܶ�<���<�1�<s�<ɰ�<���<�<)*�<3�<)*�<�<���<ɰ�<s�<�1�<���<ܶ�<��<�_�<�G�<`   `   6'�<(/�<�F�<l�<g��<���<+�<�W�<Ĕ�<���<���<��<��<��<���<���<Ĕ�<�W�<+�<���<g��<l�<�F�<(/�<`   `   �<��<�-�<;R�<��<���<{��<7�<]r�<���<���<V��<��<V��<���<���<]r�<7�<{��<���<��<;R�<�-�<��<`   `   g��<� �<��<�9�<.g�<���<���<>�<�L�<�}�<���<���<��<���<���<�}�<�L�<>�<���<���<.g�<�9�<��<� �<`   `   ���<���<"�<$�<'O�<���<9��<���<n%�<�S�<w�<��<��<��<w�<�S�<n%�<���<9��<���<'O�<$�<"�<���<`   `   ���<-��<���<R�<<;�<�i�<��<@��<J��<�)�<4J�<�^�<Df�<�^�<4J�<�)�<J��<@��<��<�i�<<;�<R�<���<-��<`   `   1��<���<\��<���<j��<�(�<�e�<���<���<Z�<�7�<DP�< Y�<DP�<�7�<Z�<���<���<�e�<�(�<j��<���<\��<���<`   `   Æ�<��<
��<��<���<��<�M�<P��<?��<��<V�<��<E!�<��<V�<��<?��<P��<�M�<��<���<��<
��<��<`   `   ���<ǟ�<%��<|��<���<��<$@�<�l�<���<y��<���<���<���<���<���<y��<���<�l�<$@�<��<���<|��<%��<ǟ�<`   `   ��<��<���<0��<��</�<L=�<�`�<ނ�<]��<���<���<���<���<���<]��<ނ�<�`�<L=�</�<��<0��<���<��<`   `   L��<���<U��<� �<&�<,�<PE�<_�<Ax�<͍�<��<��<���<��<��<͍�<Ax�<_�<PE�<,�<&�<� �<U��<���<`   `   ��<^!�<^&�<�.�<_:�<8H�<tW�<�g�<�w�<��<���<&��<���<&��<���<��<�w�<�g�<tW�<8H�<_:�<�.�<]&�<^!�<`   `   �c�<�c�<.e�<ug�<�j�<an�<Hs�<y�<�<���<��<��<ǌ�<��<��<���<�<y�<Hs�<an�<�j�<ug�<.e�<�c�<`   `   o��<̯�<���<��<��<���<���<D��<��<a��<���<��<d��<��<���<a��<��<D��<���<���<~��<��<���<̯�<`   `   ��<��<^��<���<��<���<���<ʮ�<���<t��<���<���<y��<���<���<t��<���<ʮ�<���<���<��<���<^��<��<`   `   fZ�<'V�<XJ�<�7�<u �<|�<r��<���<k��<���<w��<"��<���<"��<w��<���<k��<���<r��<|�<u �<�7�<XJ�<'V�<`   `   ���<(��<���<��<�_�<�:�<��<��<��<��<���<>��<1��<>��<���<��<��<��<��<�:�<�_�<��<���<(��<`   `   ���< ��<���<E��<��<l�<�:�<�
�<���< ��<��<���<���<���<��< ��<���<�
�<�:�<l�<��<E��<���< ��<`   `   G�<?�<�&�<� �<��<U��<J\�<W"�<T��<n��<D��<���<��<���<D��<n��<T��<W"�<J\�<U��<��<� �<�&�<?�<`   `   Ղ�<Ry�<�]�<�1�<���<��<u�<�2�<���<J��<ٝ�<,��<�~�<,��<ٝ�<J��<���<�2�<u�<��<���<�1�<�]�<Ry�<`   `   :��<x��<~��<�T�<B�<���<���<�:�<���<��<���<z�<yq�<z�<���<��<���<�:�<���<���<B�<�T�<~��<x��<`   `   ���<\��<)��<i�<�%�<U��<R��<R8�<���<̲�<��<h�<@^�<h�<��<̲�<���<R8�<R��<U��<�%�<i�<)��<\��<`   `   C��<���<ţ�<�l�<�%�<���<B�<�+�<���<���<�n�<�P�<�F�<�P�<�n�<���<���<�+�<B�<���<�%�<�l�<ţ�<���<`   `   Y��<4��<Z��<h`�<��<q��<Kl�<D�<���<���<�S�<�4�<^*�<�4�<�S�<���<���<D�<Kl�<q��<��<h`�<Z��<4��<`   `   J��<آ�<�~�<xE�<3��<y��<�O�<-��<���<g�<w4�<��<V
�<��<w4�<g�<���<-��<�O�<y��<3��<xE�<�~�<آ�<`   `   ���<gz�<�V�<h�<��<��<�+�<���<.��<BE�<�<���<���<���<�<BE�<.��<���<�+�<��<��<h�<�V�<gz�<`   `   �R�<�F�<v$�<���<���<W�<��<:��<�b�<�"�<��<���<���<���<��<�"�<�b�<:��<��<W�<���<���<v$�<�F�<`   `   u�<]�<���<���<�s�<�'�<2��<��<�?�<�<���<��<���<��<���<�<�?�<��<2��<�'�<�s�<���<���<]�<`   `   ���<��<^��<'}�<�>�<���<J��<%b�<�<_��<��<p��<.��<p��<��<_��<�<%b�<J��<���<�>�<'}�<^��<��<`   `   ���<���<�p�<�D�<��<���<���<�A�<�<���<���<��<���<��<���<���<�<�A�<���<���<��<�D�<�p�<���<`   `    Y�<DP�<�7�<Z�<���<���<�e�<�(�<j��<���<[��<���<1��<���<[��<���<j��<�(�<�e�<���<���<Z�<�7�<DP�<`   `   E!�<��<U�<��<?��<P��<�M�<��<���<��<
��<��<Æ�<��<
��<��<���<��<�M�<P��<?��<��<U�<��<`   `   ���<���<���<y��<���<�l�<$@�<��<���<|��<$��<Ɵ�<���<Ɵ�<$��<|��<���<��<$@�<�l�<���<y��<���<���<`   `   ���<���<���<]��<ނ�<�`�<L=�</�<��</��<���<��<��<��<���</��<��</�<L=�<�`�<ނ�<]��<���<���<`   `   ���<
��<��<͍�<Ax�<_�<OE�<,�<%�<� �<U��<���<K��<���<U��<� �<%�<,�<OE�<_�<Ax�<͍�<��<
��<`   `   ���<&��<���<��<�w�<�g�<tW�<8H�<_:�<�.�<]&�<]!�<��<]!�<]&�<�.�<_:�<8H�<tW�<�g�<�w�<��<���<&��<`   `   ǌ�<��<��<���<�<y�<Hs�<an�<�j�<ug�<.e�<�c�<�c�<�c�<.e�<ug�<�j�<an�<Hs�<y�<�<���<��<��<`   `   d��<��<���<a��<��<D��<���<���<~��<��<���<˯�<o��<˯�<���<��<~��<���<���<D��<��<`��<���<��<`   `   y��<���<���<t��<���<ʮ�<���<���<��<���<^��<��<��<��<^��<���<��<���<���<ʮ�<���<t��<���<���<`   `   ���<!��<w��<���<k��<���<r��<|�<u �<�7�<XJ�<'V�<fZ�<'V�<XJ�<�7�<u �<|�<r��<���<k��<���<w��<!��<`   `   1��<>��<���<��<��<��<��<�:�<�_�<��<���<(��<���<(��<���<��<�_�<�:�<��<��<��<��<���<>��<`   `   ���<���<��< ��<���<�
�<�:�<l�<��<E��<���< ��<���< ��<���<E��<��<l�<�:�<�
�<���< ��<��<���<`   `   ��<���<D��<n��<T��<W"�<J\�<U��<��<� �<�&�<?�<G�<?�<�&�<� �<��<U��<J\�<W"�<T��<n��<D��<���<`   `   �~�<,��<ٝ�<J��<���<�2�<u�<��<���<�1�<�]�<Ry�<Ղ�<Ry�<�]�<�1�<���<��<u�<�2�<���<J��<ٝ�<,��<`   `   yq�<z�<���<��<���<�:�<���<���<B�<�T�<~��<x��<:��<x��<~��<�T�<B�<���<���<�:�<���<��<���<z�<`   `   @^�<h�<��<̲�<���<R8�<S��<U��<�%�<i�<)��<\��<���<\��<)��<i�<�%�<U��<S��<R8�<���<̲�<��<h�<`   `   �F�<�P�<�n�<���<���<�+�<B�<���<�%�<�l�<ţ�<���<C��<���<ţ�<�l�<�%�<���<B�<�+�<���<���<�n�<�P�<`   `   ^*�<�4�<�S�<���<���<E�<Ll�<q��<��<h`�<Z��<4��<Y��<4��<Z��<h`�<��<q��<Ll�<D�<���<���<�S�<�4�<`   `   W
�<��<x4�<g�<���<-��<�O�<y��<3��<xE�<�~�<آ�<J��<آ�<�~�<xE�<3��<y��<�O�<-��<���<g�<x4�<��<`   `   ���<���<�<BE�<.��<���<�+�<��<��<h�<�V�<gz�<���<gz�<�V�<h�<��<��<�+�<���<.��<BE�<�<���<`   `   ���<���<��<�"�<�b�<:��<��<W�<���<���<w$�<�F�<�R�<�F�<w$�<���<���<W�<��<:��<�b�<�"�<��<���<`   `   ���<��<���<�<�?�<��<2��<�'�<�s�<���<���<]�<u�<]�<���<���<�s�<�'�<2��<��<�?�<�<���<��<`   `   .��<p��<��<_��<�<%b�<J��<���<�>�<(}�<_��<��<���<��<_��<(}�<�>�<���<J��<%b�<�<_��<��<p��<`   `   ���<��<���<���<�<�A�<���<���<��<�D�<�p�<���<���<���<�p�<�D�<��<���<���<�A�<�<���<���<��<`   `   ��<�<�2�<b�<T��<��<�:�<��<t��<��<DU�<Tw�<c��<Tw�<DU�<��<t��<��<�:�<��<T��<b�<�2�<�<`   `   ��<��<�5�<�^�<'��<���<x�<�b�<��<'��<��<�.�<V8�<�.�<��<'��<��<�b�<x�<���<'��<�^�<�5�<��<`   `   �+�<x3�<LH�<k�<���<��<d	�<RE�<_~�<!��<W��<��<u��<��<W��<!��<_~�<RE�<d	�<��<���<k�<LH�<x3�<`   `   cV�<\�<�l�<0��<���<q��<x�<!5�<	c�<���<���<��<���<��<���<���<	c�<!5�<x�<q��<���<0��<�l�<\�<`   `   {��<Y��<���<X��<��<f��<��<!4�<�U�<t�<���<��<���<��<���<t�<�U�<!4�<��<f��<��<X��<���<Y��<`   `   ^��<���<���<+��<��<K�<.)�<�?�<�T�<Ah�<Ow�<���<Ԅ�<���<Ow�<Ah�<�T�<�?�<.)�<K�<��<+��<���<���<`   `   �8�<*9�<;�<2=�<�A�<SG�<N�<�V�<C_�<�g�<�n�<s�<Tt�<s�<�n�<�g�<C_�<�V�<N�<SG�<�A�<2=�<;�<*9�<`   `   ��<���<h��<���<G��<Є�<n}�<x�<�s�<@p�<On�<]m�<yl�<]m�<On�<@p�<�s�<x�<n}�<Є�<G��<���<h��<���<`   `   ��<��<��<���<���<��<1��<7��<ӌ�<S~�<�s�<Mm�<�j�<Mm�<�s�<S~�<ӌ�<7��<1��<��<���<���<��<��<`   `   n��<�~�<�n�<�U�<w5�<b�<���<h��<r��<��<�|�<�p�<�l�<�p�<�|�<��<r��<h��<���<b�<w5�<�U�<�n�<�~�<`   `   ���<���<<��<J��<��<zY�<&�<���<���<��<م�<�t�<o�<�t�<م�<��<���<���<&�<zY�<��<J��<<��<���<`   `   �e�<�\�<@�<�<J��<���<�Z�<b�<���<@��<��<�u�<�n�<�u�<��<@��<���<b�<�Z�<���<J��<�<@�<�\�<`   `   3��<��<ؚ�<�f�<|#�<,��<ˆ�<�9�<���<:��<�<�r�<�i�<�r�<�<:��<���<�9�<ˆ�<,��<|#�<�f�<ؚ�<��<`   `   �<��<���<b��<5\�<��<e��<�O�<���<A��<��<;i�<*^�<;i�<��<A��<���<�O�<e��<��<5\�<b��<���<��<`   `   ^W�<�H�<��<!��<a��<#�<���<1Y�<���<���<~{�<MX�<GL�<MX�<~{�<���<���<1Y�<���<#�<a��<!��<��<�H�<`   `   �|�< m�<�>�<���<*��<�/�<��<�U�<��<ˢ�<ae�<�?�<+3�<�?�<ae�<ˢ�<��<�U�<��<�/�<*��<���<�>�< m�<`   `   P��<#x�<�G�<��<���<R*�<N��<nE�<���<ƈ�<�G�<��<g�<��<�G�<ƈ�<���<nE�<N��<R*�<���<��<�G�<#x�<`   `   �{�<�j�<�8�<���<���<.�<��<�(�<k��<�e�<|#�<��<��<��<|#�<�e�<k��<�(�<��<.�<���<���<�8�<�j�<`   `   X�<zF�<`�<���<a�<<��<�u�<� �<L��<�<�<���<���<���<���<���<�<�<L��<� �<�u�<<��<a�<���<`�<zF�<`   `   ��<Q�<5��<��<{,�<|��<�D�<��<Vh�<�<)��<��<��<��<)��<�<Uh�<��<�D�<|��<{,�<��<5��<Q�<`   `   ��<���<���<M�<Q��<��<3�<G��<�7�<���<E��<Yy�<�k�<Yy�<E��<���<�7�<G��<3�<��<Q��<M�<���<���<`   `   ���<u�<]H�<��<I��<b?�<���<�h�<��<ݵ�<�x�<lR�<E�<lR�<�x�<ݵ�<��<�h�<���<b?�<I��<��<]H�<u�<`   `   -�<I�<d��<i��<�_�<��<���<7�<=��<C��<@W�<3�<'�<3�<@W�<C��<=��<7�<���<��<�_�<i��<d��<I�<`   `   ���<���<Ϣ�<�f�<g�<���<Wf�<��<θ�<�s�<�>�<��<��<��<�>�<�s�<θ�<��<Wf�<���<g�<�f�<Ϣ�<���<`   `   b��<Tw�<DU�<��<t��<��<�:�<��<S��<b�<�2�<�<��<�<�2�<b�<S��<��<�:�<��<t��<��<DU�<Tw�<`   `   V8�<�.�<��<'��<��<�b�<x�<���<&��<�^�<�5�<��<��<��<�5�<�^�<&��<���<x�<�b�<��<'��<��<�.�<`   `   u��<��<W��<!��<_~�<RE�<d	�<��<���<k�<LH�<x3�<�+�<x3�<LH�<k�<���<��<d	�<RE�<_~�<!��<W��<��<`   `   ���<��<���<���<	c�<!5�<x�<p��<���</��<�l�<\�<cV�<\�<�l�</��<���<p��<x�<!5�<	c�<���<���<��<`   `   ���<��<���<t�<�U�<!4�<��<f��<��<X��<���<X��<{��<X��<���<X��<��<f��<��<!4�<�U�<t�<���<��<`   `   Ԅ�<���<Ow�<Ah�<�T�<�?�<.)�<K�<��<+��<���<���<^��<���<���<+��<��<K�<.)�<�?�<�T�<Ah�<Ow�<���<`   `   Tt�<s�<�n�<�g�<C_�<�V�<N�<SG�<�A�<2=�<;�<*9�<�8�<*9�<;�<2=�<�A�<SG�<N�<�V�<C_�<�g�<�n�<s�<`   `   yl�<]m�<On�<@p�<�s�<x�<n}�<Є�<G��<���<h��<���<��<���<h��<���<G��<Є�<n}�<x�<�s�<@p�<On�<]m�<`   `   �j�<Lm�<�s�<S~�<ӌ�<7��<1��<��<���<���<��<��<��<��<��<���<���<��<1��<7��<ӌ�<S~�<�s�<Lm�<`   `   �l�<�p�<�|�<��<r��<h��<���<b�<w5�<�U�<�n�<�~�<n��<�~�<�n�<�U�<w5�<b�<���<h��<r��<��<�|�<�p�<`   `   o�<�t�<؅�<��<���<���<&�<zY�<��<J��<<��<���<���<���<<��<J��<��<zY�<&�<���<���<��<؅�<�t�<`   `   �n�<�u�<��<@��<���<b�<�Z�<���<J��<�<@�<�\�<�e�<�\�<@�<�<J��<���<�Z�<b�<���<@��<��<�u�<`   `   �i�<�r�<�<:��<���<�9�<ˆ�<,��<|#�<�f�<ؚ�<��<3��<��<ؚ�<�f�<|#�<,��<ˆ�<�9�<���<:��<�<�r�<`   `   *^�<;i�<��<A��<���<�O�<e��<��<5\�<c��<���<��<�<��<���<c��<5\�<��<e��<�O�<���<A��<��<;i�<`   `   GL�<MX�<~{�<���<���<1Y�<���<#�<a��<!��<��<�H�<^W�<�H�<��<!��<a��<#�<���<1Y�<���<���<~{�<MX�<`   `   +3�<�?�<ae�<ˢ�<��<�U�<��<�/�<*��<���<�>�< m�<�|�< m�<�>�<���<*��<�/�<��<�U�<��<ˢ�<ae�<�?�<`   `   g�<��<�G�<ƈ�<���<nE�<O��<R*�<���<��<�G�<#x�<P��<#x�<�G�<��<���<R*�<O��<nE�<���<ƈ�<�G�<��<`   `   ��<��<|#�<�e�<k��<�(�<��<.�<���<���<�8�<�j�<�{�<�j�<�8�<���<���<.�<��<�(�<k��<�e�<|#�<��<`   `   ���<���<���<�<�<L��<� �<�u�<=��<a�<���<`�<{F�<X�<{F�<`�<���<a�<=��<�u�<� �<L��<�<�<���<���<`   `   ��<��<)��<�<Vh�<��<�D�<|��<{,�<��<5��<Q�<��<Q�<5��<��<{,�<|��<�D�<��<Vh�<�<)��<��<`   `   �k�<Yy�<E��<���<�7�<G��<3�<��<Q��<M�<���<���<��<���<���<M�<Q��<��<3�<G��<�7�<���<E��<Yy�<`   `   E�<lR�<�x�<ݵ�<��<�h�<���<b?�<I��<��<]H�<u�<���<u�<]H�<��<I��<b?�<���<�h�<��<ݵ�<�x�<lR�<`   `   '�<3�<@W�<C��<=��<7�<���<��<�_�<i��<d��<I�<-�<I�<d��<i��<�_�<��<���<7�<=��<C��<@W�<3�<`   `   ��<��<�>�<�s�<θ�<��<Wf�<���<g�<�f�<Ϣ�<���<���<���<Ϣ�<�f�<g�<���<Wf�<��<θ�<�s�<�>�<��<`   `   o�<�{�<G��<���<2�<���<���<hm�<���<3�<�z�<̨�<���<̨�<�z�<3�<���<hm�<���<���<2�<���<G��<�{�<`   `   y�<���<���<���<Z#�<1x�<H��<!5�<���<���<��<=F�<�S�<=F�<��<���<���<!5�<H��<1x�<Z#�<���<���<���<`   `   ��<���<[��<���<�'�<�o�<���<5�<[�<)��<���<���<��<���<���<)��<[�<5�<���<�o�<�'�<���<[��<���<`   `   ���<���<��<��<7A�<�z�<ݸ�<���<�7�<m�<��<��<��<��<��<m�<�7�<���<ݸ�<�z�<7A�<��<��<���<`   `   r�<�#�<�3�<N�<�p�<��<���<���<&&�<]N�<�n�<���<T��<���<�n�<]N�<&&�<���<���<��<�p�<N�<�3�<�#�<`   `   ���<��<M��<k��<j��<���<���<[�<�%�<T@�<�U�<c�<Ng�<c�<�U�<T@�<�%�<[�<���<���<j��<k��<M��<��<`   `   ���<n��<s��<6�<a�<��<��<�'�<Z4�<�@�<mJ�<�Q�<�S�<�Q�<mJ�<�@�<Z4�<�'�<��<��<a�<6�<s��<n��<`   `   ���<Ѓ�<k~�<-v�<�l�<�b�<:Z�<�R�<�N�<DL�<�J�<�J�< K�<�J�<�J�<DL�<�N�<�R�<:Z�<�b�<�l�<-v�<k~�<Ѓ�<`   `   �<F�<N
�<��<b��<��<-��<���<Pq�<�_�<�R�<�K�<YI�<�K�<�R�<�_�<Pq�<���<-��<��<b��<��<N
�<F�<`   `   ��<$��<Ȝ�<�z�<�O�<
 �<���<���<��<mv�<E^�<�O�<�J�<�O�<E^�<mv�<��<���<���<
 �<�O�<�z�<Ȝ�<$��<`   `   ZX�<�M�<�/�<d �<���<I��<�:�<���<"��<��<hi�<�S�<�K�<�S�<hi�<��<"��<���<�:�<I��<���<d �<�/�<�M�<`   `   ���<C��<���<�~�<�1�<(��<ہ�<�+�<���<f��<kq�<�T�<OJ�<�T�<kq�<f��<���<�+�<ہ�<(��<�1�<�~�<���<C��<`   `   kv�<Rf�<�7�<���<���<A*�<O��<(V�<���<$��<�r�<fO�<TC�<fO�<�r�<$��<���<(V�<O��<A*�<���<���<�7�<Rf�<`   `   o��<���<ٟ�<�K�<��<�h�<���<s�<��<<��<j�<.A�<93�<.A�<j�<<��<��<s�<���<�h�<��<�K�<ٟ�<���<`   `   �;�<0'�<d��<^��<X�<��<��<��<w�<ݢ�<zW�<�)�<��<�)�<zW�<ݢ�<w�<��<��<��<X�<^��<d��<0'�<`   `   �p�<�Y�<��<e��<5�<ѣ�<1�<�{�<���<���<-:�<S�<-��<S�<-:�<���<���<�{�<1�<ѣ�<5�<e��<��<�Y�<`   `   ���<Ij�<2&�<���<6�<6��<���<e�<���<�g�<��<���<V��<���<��<�g�<���<e�<���<6��<6�<���<2&�<Ij�<`   `   jo�<zW�<�<ԥ�<v�<�~�<]��<:=�<:��<�8�<D��<w��<���<w��<D��<�8�<:��<:=�<]��<�~�<v�<ԥ�<�<zW�<`   `   z<�<�$�<���<�r�<&��<�J�<Ԧ�<�<Cy�<{�<\��<�q�<�^�<�q�<\��<{�<Cy�<�<Ԧ�<�J�<&��<�r�<���<�$�<`   `   ���<=��<>��<](�<%��<��<�d�<s��<S;�<x��<�m�</7�<B$�</7�<�m�<x��<S;�<s��<�d�<��<%��<](�<>��<=��<`   `   6��<�t�<�2�<@��<5I�<���<��<W��<0��<܈�<A3�<|��<���<|��<A3�<܈�<0��<W��<��<���<5I�<@��<�2�<�t�<`   `   2�<��<��<�e�<���<K]�<}��<�;�<���<�N�<��<���<i��<���<��<�N�<���<�;�<}��<K]�<���<�e�<��<��<`   `   ���<Ԍ�<�S�<���<��<��<�}�<F��<&��<�<���<���<@��<���<���<�<&��<F��<�}�<��<��<���<�S�<Ԍ�<`   `   �(�<0�<P��<d��<U*�<A��<u8�<��<�R�<���<��<{��<Lx�<{��<��<���<�R�<��<u8�<A��<U*�<d��<P��<0�<`   `   ���<̨�<�z�<3�<���<hm�<���<���<2�<���<G��<�{�<o�<�{�<G��<���<2�<���<���<hm�<���<3�<�z�<̨�<`   `   �S�<<F�<��<���<���<!5�<H��<0x�<Z#�<���<���<���<y�<���<���<���<Z#�<0x�<H��<!5�<���<���<��<<F�<`   `   ��<���<���<)��<[�<5�<���<�o�<�'�<���<[��<���<��<���<[��<���<�'�<�o�<���<5�<[�<)��<���<���<`   `   ��<��<��<m�<�7�<���<ݸ�<�z�<7A�<��<��<���<���<���<��<��<7A�<�z�<ݸ�<���<�7�<m�<��<��<`   `   S��<���<�n�<]N�<&&�<���<���<��<�p�<N�<�3�<�#�<r�<�#�<�3�<N�<�p�<��<���<���<&&�<]N�<�n�<���<`   `   Mg�<c�<�U�<S@�<�%�<[�<���<���<i��<k��<M��<��<���<��<M��<k��<i��<���<���<[�<�%�<S@�<�U�<c�<`   `   �S�<�Q�<mJ�<�@�<Z4�<�'�<��<��<a�<6�<s��<m��<���<m��<s��<6�<a�<��<��<�'�<Z4�<�@�<mJ�<�Q�<`   `    K�<�J�<�J�<DL�<�N�<�R�<:Z�<�b�<�l�<-v�<k~�<σ�<���<σ�<k~�<-v�<�l�<�b�<:Z�<�R�<�N�<DL�<�J�<�J�<`   `   YI�<�K�<�R�<�_�<Pq�<���<,��<��<b��<��<N
�<F�<�<F�<N
�<��<b��<��<,��<���<Pq�<�_�<�R�<�K�<`   `   �J�<�O�<E^�<mv�<��<���<���<
 �<�O�<�z�<ǜ�<$��<��<$��<ǜ�<�z�<�O�<
 �<���<���<��<mv�<E^�<�O�<`   `   �K�<�S�<hi�<��<"��<���<�:�<H��<���<d �<�/�<�M�<ZX�<�M�<�/�<d �<���<H��<�:�<���<"��<��<hi�<�S�<`   `   OJ�<�T�<kq�<f��<���<�+�<ہ�<(��<�1�<�~�<���<C��<���<C��<���<�~�<�1�<(��<ہ�<�+�<���<f��<kq�<�T�<`   `   TC�<fO�<�r�<$��<���<(V�<O��<A*�<���<���<�7�<Rf�<kv�<Rf�<�7�<���<���<A*�<O��<(V�<���<$��<�r�<fO�<`   `   93�<.A�<j�<<��<��<s�<���<�h�<��<�K�<ٟ�<���<o��<���<ٟ�<�K�<��<�h�<���<s�<��<<��<j�<.A�<`   `   ��<�)�<zW�<ݢ�<w�<��<��<��<X�<^��<d��<0'�<�;�<0'�<d��<^��<X�<��<��<��<w�<ݢ�<zW�<�)�<`   `   -��<S�<-:�<���<���<�{�<1�<ѣ�<5�<e��<��<�Y�<�p�<�Y�<��<e��<5�<ѣ�<1�<�{�<���<���<-:�<S�<`   `   V��<���<��<�g�<���<e�<���<6��<6�<���<2&�<Ij�<���<Ij�<2&�<���<6�<6��<���<e�<���<�g�<��<���<`   `   ���<x��<E��<�8�<:��<:=�<^��<�~�<v�<ԥ�<�<zW�<ko�<zW�<�<ԥ�<v�<�~�<]��<:=�<:��<�8�<E��<w��<`   `   �^�<�q�<\��<{�<Cy�<�<Ԧ�<�J�<&��<�r�<���<�$�<z<�<�$�<���<�r�<&��<�J�<Ԧ�<�<Cy�<{�<\��<�q�<`   `   B$�</7�<�m�<x��<S;�<s��<�d�<��<&��<](�<?��<=��<���<=��<?��<](�<&��<��<�d�<s��<S;�<x��<�m�</7�<`   `   ���<|��<A3�<܈�<1��<W��<��<���<5I�<A��<�2�<�t�<6��<�t�<�2�<@��<5I�<���<��<W��<0��<܈�<A3�<|��<`   `   i��<���<��<�N�<���<�;�<}��<K]�<���<�e�<��<��<2�<��<��<�e�<���<K]�<}��<�;�<���<�N�<��<���<`   `   @��<���<���<�<&��<G��<�}�<��<��<���<�S�<Ԍ�<���<Ԍ�<�S�<���<��<��<�}�<G��<&��<�<���<���<`   `   Lx�<{��<��<���<�R�<��<v8�<A��<V*�<d��<P��<0�<�(�<0�<P��<d��<U*�<A��<v8�<��<�R�<���<��<{��<`   `   ���<P��<$��<I1�<��<t�<@��<�?�<��<�H�<ϩ�<���<1��<���<ϩ�<�H�<��<�?�<@��<t�<��<I1�<$��<P��<`   `   f��<9��<���<,�<���<e��<Qu�<���<-n�<f��<�.�<Hd�<�v�<Hd�<�.�<f��<-n�<���<Qu�<e��<���<,�<���<9��<`   `   5��<���<q�<�A�<K��<���<�V�<���<R(�<(��<���<��<��<��<���<(��<R(�<���<�V�<���<K��<�A�<q�<���<`   `   ��<h&�<�C�<Ds�<���<���<
R�<#��<��<�C�<�|�<���<­�<���<�|�<�C�<��<#��<
R�<���<���<Ds�<�C�<h&�<`   `   |��<��<S��<���<e��<c(�<~f�<���<c��<b�<�G�<d�<m�<d�<�G�<b�<c��<���<}f�<c(�<e��<���<S��<��<`   `   �<��<��<,�<�H�<Yk�<��<���<���<��<�(�<[<�<�B�<[<�<�(�<��<���<���<��<Yk�<�H�<,�<��<��<`   `   ߦ�<ʧ�<]��<Ȱ�<o��<D��<_��<W��<D��<0�<�<>&�<q)�<>&�<�<0�<D��<W��<_��<D��<o��<Ȱ�<]��<ʧ�<`   `   �^�<�\�<U�<K�<\>�<�1�<�(�<�!�<��<��<��<��<��<��<��<��<��<�!�<�(�<�1�<\>�<K�<U�<�\�<`   `   +)�<�#�<��<���<X��<Ǭ�<���<sg�<�K�<�6�<!(�<��<�<��<!(�<�6�<�K�<sg�<���<Ǭ�<X��<���<��<�#�<`   `   t��<���<���<���<�n�<'/�<���<��<�~�<U�<�6�<$�<0�<$�<�6�<U�<�~�<��<���<'/�<�n�<���<���<���<`   `   %��<l��<���<�]�<��<I��<�T�<���<Ȱ�<Nr�<!E�<[)�< �<[)�<!E�<Nr�<Ȱ�<���<�T�<I��<��<�]�<���<l��<`   `   N��<Y��<^�<�
�<-��<.,�<���<B�<���<u��<�M�<�(�<��<�(�<�M�<u��<���<B�<���<.,�<-��<�
�<^�<Y��<`   `   Va�<�J�<�
�<Q��<�%�<���<�<�y�<���<���<*M�<e�<k�<e�<*M�<���<���<�y�<�<���<�%�<Q��<�
�<�J�<`   `   ���<���<��<�%�<$��<���<oB�<ڟ�<]�<��<�@�<��<���<��<�@�<��<]�<ڟ�<oB�<���<$��<�%�<��<���<`   `   �v�<�Y�<��<8��<G��<)%�<�f�<���<��<Z��<�&�<4��<s��<4��<�&�<Z��<��<���<�f�<)%�<G��<8��<��<�Y�<`   `   P��<>��<�E�<��<z�<�=�<Wo�<���<���<�h�<u��<���<̤�<���<u��<�h�<���<���<Wo�<�=�<z�<��<�E�<>��<`   `   ���<r��<X�<��<.�<15�<�[�<V��<}��<�7�<���<$��<�i�<$��<���<�7�<}��<V��<�[�<15�<.�<��<X�<r��<`   `   ���<���<�;�<���<%��<=�<�+�<�U�<���<���<E��<�<�<�$�<�<�<E��<���<���<�U�<�+�<=�<%��<���<�;�<���<`   `   (w�<�U�<���<�\�<���<;��<���<�<�N�<��<�9�<w��<t��<w��<�9�<��<�N�<�<���<;��<���<�\�<���<�U�<`   `   	�<���<��<���<	:�<Ze�<a��<R��<<��<4_�<��<3��<��<3��<��<4_�<<��<R��<a��<Ze�<	:�<���<��<���<`   `   �}�<�^�<,�<Dv�<R��<���<\$�<�Z�<��<��<���<�Y�<=B�<�Y�<���<��<��<�Z�<\$�<���<R��<Dv�<,�<�^�<`   `   k��<��<�m�<���<�?�<��<��<C��<)Q�<���<#X�<�<�<�<#X�<���<)Q�<C��<��<��<�?�<���<�m�<��<`   `   �9�<W�<p��<mV�<���<�<ET�<���<@�<���<�<~��<���<~��<�<���<@�<���<ET�<�<���<mV�<p��<W�<`   `   ��<�}�<*7�<0��<�<�<���<���<�W�<���<�N�<O��<���<{��<���<O��<�N�<���<�W�<���<���<�<�<0��<*7�<�}�<`   `   1��<���<ϩ�<�H�<��<�?�<@��<s�<��<H1�<$��<P��<���<P��<$��<H1�<��<s�<@��<�?�<��<�H�<ϩ�<���<`   `   �v�<Hd�<�.�<f��<-n�<���<Pu�<e��<���<,�<���<9��<f��<9��<���<,�<���<e��<Pu�<���<-n�<f��<�.�<Hd�<`   `   ��<��<���<(��<R(�<���<�V�<���<K��<�A�<q�<���<4��<���<q�<�A�<K��<���<�V�<���<Q(�<(��<���<��<`   `   ���<���<�|�<�C�<��<"��<
R�<���<���<Ds�<�C�<h&�<��<h&�<�C�<Ds�<���<���<
R�<"��<��<�C�<�|�<���<`   `   m�<d�<�G�<b�<b��<���<}f�<c(�<e��<���<S��<��<|��<��<R��<���<d��<c(�<}f�<���<b��<b�<�G�<d�<`   `   �B�<[<�<�(�<��<���<���<��<Xk�<�H�<,�<��<��<�<��<��<,�<�H�<Xk�<��<���<���<��<�(�<Z<�<`   `   q)�<>&�<�</�<D��<W��<^��<C��<o��<Ȱ�<]��<ʧ�<ߦ�<ʧ�<]��<Ȱ�<o��<C��<^��<W��<D��</�<�<>&�<`   `   ��<��<��<��<��<�!�<�(�<�1�<\>�<K�<U�<�\�<�^�<�\�<U�<K�<\>�<�1�<�(�<�!�<��<��<��<��<`   `   �<��<!(�<�6�<�K�<sg�<���<Ǭ�<X��<���<��<�#�<+)�<�#�<��<���<X��<Ǭ�<���<sg�<�K�<�6�<!(�<��<`   `   0�<$�<�6�<U�<�~�<��<���<'/�<�n�<��<���<���<t��<���<���<��<�n�<'/�<���<��<�~�<U�<�6�<$�<`   `    �<[)�<!E�<Nr�<ǰ�<���<�T�<I��<��<�]�<���<l��<%��<l��<���<�]�<��<I��<�T�<���<ǰ�<Nr�<!E�<Z)�<`   `   ��<�(�<�M�<u��<���<B�<���<.,�<-��<�
�<^�<Y��<N��<Y��<^�<�
�<-��<.,�<���<B�<���<u��<�M�<�(�<`   `   k�<e�<*M�<���<���<�y�<�<���<�%�<Q��<�
�<�J�<Va�<�J�<�
�<Q��<�%�<���<�<�y�<���<���<*M�<e�<`   `   ���<��<�@�<��<]�<ڟ�<oB�<���<$��<�%�<��<���<���<���<��<�%�<$��<���<oB�<ڟ�<]�<��<�@�<��<`   `   s��<4��<�&�<Z��<��<���<�f�<)%�<G��<8��<��<�Y�<�v�<�Y�<��<8��<G��<)%�<�f�<���<��<Z��<�&�<4��<`   `   ͤ�<���<u��<�h�<���< ��<Wo�<�=�<z�<��<�E�<>��<P��<>��<�E�<��<z�<�=�<Wo�<���<���<�h�<u��<���<`   `   �i�<$��<���<�7�<}��<V��<�[�<15�<.�<��<X�<r��<���<r��<X�<��<.�<15�<�[�<V��<}��<�7�<���<$��<`   `   �$�<�<�<E��<���<���<�U�<�+�<=�<%��<���<�;�<���<���<���<�;�<���<%��<=�<�+�<�U�<���<���<E��<�<�<`   `   t��<x��<�9�<��<�N�<�<���<;��<���<�\�<���<�U�<(w�<�U�<���<�\�<���<;��<���<�<�N�<��<�9�<x��<`   `   ��<4��<��<4_�<<��<R��<a��<Ze�<	:�<���<��<���<	�<���<��<���<	:�<Ze�<a��<R��<<��<4_�<��<4��<`   `   =B�<�Y�<���<��<��<�Z�<\$�<���<R��<Ev�<,�<�^�<�}�<�^�<,�<Ev�<R��<���<\$�<�Z�<��<��<���<�Y�<`   `   �<�<#X�<���<*Q�<D��<��<��<�?�<���<�m�<��<k��<��<�m�<���<�?�<��<��<D��<*Q�<���<#X�<�<`   `   ���<~��<�<���<@�<���<ET�<�<���<nV�<p��<W�<�9�<W�<p��<nV�<���<�<ET�<���<@�<���<�<~��<`   `   {��<���<O��<�N�<���<�W�<���<���<�<�<0��<*7�<�}�<��<�}�<*7�<0��<�<�<���<���<�W�<���<�N�<O��<���<`   `   ��<���<���<�H�<#��<�|�<d8�<��<P��<n_�<i��<�7�<T�<�7�<i��<n_�<P��<��<d8�<�|�<#��<�H�<���<���<`   `   ���<���<���<�A�<߻�<xN�<k��<v��<w=�<���<�>�<���<���<���<�>�<���<w=�<v��<j��<xN�<߻�<�A�<���<���<`   `   g��<j��<��<^�<M��<�@�<d��<DY�<^��<�[�<3��<'��<9�<'��<3��<�[�<^��<DY�<d��<�@�<M��<^�<��<j��<`   `   -�<_:�<�`�<��<!��<pU�<���<�8�<ڧ�<�
�<-W�<l��<k��<l��<-W�<�
�<ڧ�<�8�<���<pU�<!��<��<�`�<_:�<`   `   ��<��<��<-�<�B�<|��<w��<k9�<��<���<Y�<R:�<�G�<R:�<Y�<���<��<k9�<w��<|��<�B�<-�<��<��<`   `   @]�<1c�<ct�<���<��<���<��<�W�<<��<��<��<��<)�<��<��<��<<��<�W�<��<���<��<���<ct�<1c�<`   `   z/�<1�<�5�<=>�<DK�<7^�<u�<���<N��<t��<���<���<���<���<���<t��<N��<���<u�<7^�<DK�<=>�<�5�<1�<`   `   �$�<!�<j�<�	�<���<A��<���<���<I��<���<���<^��<���<^��<���<���<I��<���<���<A��<���<�	�<j�<!�<`   `   m4�<,�<L�<!��<���<ʐ�<�b�<n:�<��<�<V��<���<���<���<V��<�<��<n:�<�b�<ʐ�<���<!��<L�<,�<`   `   JV�<~H�<��<��<��<#>�<)��<��<�[�<z(�<��<h��<��<h��<��<z(�<�[�<��<)��<#>�<��<��<��<~H�<`   `   �|�<j�<0�<���<�g�<���<�r�<. �<	��<[N�<U�<���<���<���<U�<[N�<	��<. �<�r�<���<�g�<���<0�<j�<`   `   ���<�|�<22�<!��<�3�<ȓ�<���<�Z�<'��<�k�<��<���<���<���<��<�k�<'��<�Z�<���<ȓ�<�3�<!��<22�<�|�<`   `   ���<�|�<�!�<f��<]��<�%�<x^�<1��<\ �<�{�<��<���<@��<���<��<�{�<\ �<1��<x^�<�%�<]��<f��<�!�<�|�<`   `   �x�<HT�<���<�G�<Wz�<T��<ܱ�<���<Z�<gz�<��<���<«�<���<��<gz�<Z�<���<ܱ�<T��<Wz�<�G�<���<HT�<`   `   ��<t��<k��<���<���<:��<��<
��<��<�c�<���<|��<-z�<|��<���<�c�<��<
��<��<:��<���<���<k��<t��<`   `   E��<�[�<'��<��<H�</�<}��<��<���<	7�<��<*T�<�7�<*T�<��<	7�<���<��<}��</�<H�<��<'��<�[�<`   `   8��<2{�<���<�$�<��<O��<���<W��<���<���<�_�<��<���<��<�_�<���<���<W��<���<O��<��<�$�<���<2{�<`   `   ���<LV�<��<���<���<Y��<[��<2q�<Op�<4��<6�<=��<���<=��<6�<4��<Op�<2q�<[��<Y��<���<���<��<LV�<`   `   �!�<H��<�i�<��<��<:d�<52�<N�<9�<=�<��<mD�<	%�<mD�<��<=�<9�<N�<52�<:d�<��<��<�i�<H��<`   `   ���<�X�<���<��<�<���<ѷ�<˛�<_��<��<\;�<���<C��<���<\;�<��<_��<˛�<ѷ�<���<�<��<���<�X�<`   `   ��<n��<$�<JT�<�a�<lK�<�-�<v�<f-�<�g�<H��<`}�<q_�<`}�<H��<�g�<f-�<v�<�-�<lK�<�a�<JT�<$�<n��<`   `   ��<n��<�G�<���<B��<s��<5��<[��<ս�<�<�z�<�&�<�	�<�&�<�z�<�<ս�<[��<5��<s��<B��<���<�G�<n��<`   `   n�<��<�t�<���<W��<�
�<�<�+�<�Z�<���<�.�<���<��<���<�.�<���<�Z�<�+�<�<�
�<W��<���<�t�<��<`   `   6#�<��<���<��<�N�<x�<ț�<��<�
�<>n�<���<���<~��<���<���<>n�<�
�<��<ț�<x�<�N�<��<���<��<`   `   T�<�7�<i��<n_�<P��<��<d8�<�|�<#��<�H�<���<���<��<���<���<�H�<"��<�|�<d8�<��<P��<n_�<i��<�7�<`   `   ���<���<�>�<���<w=�<v��<j��<wN�<޻�<�A�<���<���<���<���<���<�A�<޻�<wN�<j��<v��<w=�<���<�>�<���<`   `   9�<&��<3��<�[�<^��<DY�<c��<�@�<L��<^�<��<j��<f��<j��<��<^�<L��<�@�<c��<CY�<]��<�[�<3��<&��<`   `   k��<l��<-W�<�
�<٧�<�8�<���<pU�<!��<��<�`�<_:�<-�<_:�<�`�<��<!��<pU�<���<�8�<٧�<�
�<-W�<l��<`   `   �G�<R:�<X�<���<��<k9�<w��<{��<�B�<,�<��<��<��<��<��<,�<�B�<{��<w��<k9�<��<���<X�<R:�<`   `   (�<��<��<��<<��<�W�<��<���<��<���<ct�<1c�<@]�<1c�<ct�<���<��<���<��<�W�<<��<��<��<��<`   `   ���<���<���<t��<N��<���<u�<6^�<DK�<=>�<�5�<1�<z/�<1�<�5�<=>�<DK�<6^�<u�<���<N��<t��<���<���<`   `   ���<^��<���<���<I��<���<���<A��<���<�	�<i�<!�<�$�<!�<i�<�	�<���<A��<���<���<I��<���<���<^��<`   `   ���<���<U��<�<��<n:�<�b�<ʐ�<���<!��<L�<,�<m4�<,�<L�<!��<���<ʐ�<�b�<n:�<��<�<U��<���<`   `   ��<h��<��<z(�<�[�<��<)��<#>�<��<��<��<~H�<IV�<~H�<��<��<��<">�<)��<��<�[�<z(�<��<h��<`   `   ���<���<U�<[N�<	��<. �<�r�<���<�g�<���<0�<j�<�|�<j�<0�<���<�g�<���<�r�<. �<	��<[N�<U�<���<`   `   ���<���<��<�k�<'��<�Z�<���<ȓ�<�3�<!��<22�<�|�<���<�|�<22�<!��<�3�<ȓ�<���<�Z�<'��<�k�<��<���<`   `   @��<���<��<�{�<\ �<1��<x^�<�%�<]��<f��<�!�<�|�<���<�|�<�!�<f��<]��<�%�<x^�<1��<\ �<�{�<��<���<`   `   «�<���<��<gz�<Z�<���<ܱ�<T��<Xz�<�G�<���<IT�<�x�<HT�<���<�G�<Wz�<T��<ܱ�<���<Z�<gz�<��<���<`   `   -z�<|��<���<�c�<��<
��<��<:��<���<���<k��<t��<��<t��<k��<���<���<:��<��<
��<��<�c�<���<|��<`   `   �7�<*T�<��<	7�<���<��<}��<0�<H�<��<(��<�[�<E��<�[�<(��<��<H�</�<}��<��<���<	7�<��<*T�<`   `   ���<��<�_�<���<���<W��<���<O��<��<�$�<���<2{�<8��<2{�<���<�$�<��<O��<���<W��<���<���<�_�<��<`   `   ���<>��<6�<4��<Op�<2q�<\��<Z��<���<���<��<LV�<���<LV�<��<���<���<Z��<\��<2q�<Op�<4��<6�<>��<`   `   	%�<mD�<��<=�<9�<N�<52�<:d�<���<��<�i�<I��<�!�<I��<�i�<��<���<:d�<52�<N�<9�<=�<��<mD�<`   `   C��<���<];�<��<_��<˛�<ҷ�<���<�<��<���<�X�<���<�X�<���<��<�<���<ѷ�<˛�<_��<��<];�<���<`   `   q_�<a}�<H��<�g�<f-�<v�<�-�<lK�<�a�<JT�<%�<o��<��<o��<%�<JT�<�a�<lK�<�-�<v�<f-�<�g�<H��<a}�<`   `   �	�<�&�<�z�<�<ս�<[��<6��<s��<C��<���<�G�<n��<��<n��<�G�<���<C��<s��<5��<[��<ս�<�<�z�<�&�<`   `   ��<���<�.�<���<�Z�<�+�<�<�
�<W��<���<�t�<��<o�<��<�t�<���<W��<�
�<�<�+�<�Z�<���<�.�<���<`   `   ~��<���<���<?n�<�
�<��<ț�<x�<�N�<��<���<��<7#�<��<���<��<�N�<x�<ț�<��<�
�<?n�<���<���<`   `   � �<�<�<ڍ�<��<h��<[��<ݖ�<��<��<�p�<|"�<��<Ǽ�<��<|"�<�p�<��<��<ݖ�<[��<h��<��<ڍ�<�<�<`   `   �6�<{O�<��<�<&��<�f�<M<�<~�<���<i��<�I�<���<���<���<�I�<i��<���<~�<M<�<�f�<&��<�<��<{O�<`   `   �y�<R��<y��<�/�<:��<�X�<��<��<G�<� �<��<���<c�<���<��<� �<G�<��<��<�X�<:��<�/�<y��<R��<`   `   ���<. �<+2�<���<���<v�<?	�<q��<�6�<C��<�"�<ze�<'|�<ze�<�"�<C��<�6�<q��<?	�<v�<���<���<+2�<. �<`   `   ���<���<���<��<K[�<��<�0�<���<L�<H�<<��<��<��<��<<��<H�<L�<���<�0�<��<K[�<��<���<���<`   `   <v�<L}�<��<%��<���<84�<��<���<e!�<�i�<���<&��<G��<&��<���<�i�<e!�<���<��<84�<���<%��<��<L}�<`   `   ���<���<C��<מ�<��<���<���<��<yH�<Mr�<Ô�<Ȫ�<v��<Ȫ�<Ô�<Lr�<yH�<��<���<���<��<מ�<C��<���<`   `   ���<:��<k��<̫�<���<��<���<���<+��<Q��<͚�<��<\��<��<͚�<Q��<+��<���<���<��<���<̫�<j��<:��<`   `   w2�<�&�<'�<���<1��<�c�<�*�<���<4��<ʽ�<��<إ�<&��<إ�<��<ʽ�<4��<���<�*�<�c�<1��<���<'�<�&�<`   `   ���<O��<p�<�<���<zE�<���<)}�<"-�<���< ��<έ�<��<έ�< ��<���<"-�<)}�<���<zE�<���<�<p�<O��<`   `   �L�<�1�<��<j�<��<
0�<q��<���<@��<��<D��<Q��<S��<Q��<D��<��<@��<���<q��<
0�<��<j�<��<�1�<`   `   ���<���<�K�<��<��<U�<�7�<�t�<���<�B�<���<Ǩ�<ە�<Ǩ�<���<�B�<���<�t�<�7�<U�<��<��<�K�<���<`   `   �<�<��<���<���<���<���<��<���<I��<\T�<���<��<�x�<��<���<\T�<H��<���<��<���<���<���<���<��<`   `   �l�<�:�<ҩ�<���<9��<�u�<:�<��<��<N�<���<1d�<�F�<0d�<���<N�<��<��<:�<�u�<9��<���<ҩ�<�:�<`   `   ?R�<��<�x�<{}�<0@�<G��<9|�<�.�<��<I,�<Q��<�!�<� �<�!�<Q��<I,�<��<�.�<9|�<G��<0@�<{}�<�x�<��<`   `   ���<"��<���<���<��<7�<��<� �<��<��<�6�<0��<���<0��<�6�<��<��<� �<��<7�<��<���<���<"��<`   `   ��<���<}�<e��<0��<N��<f�<"��<���<���<���<]�<�6�<]�<���<���<���<"��<f�<N��<0��<e��<}�<���<`   `   C��<D��<9��<���<"K�<���<{�<<��<�0�<� �<�Y�<��<߹�<��<�Y�<� �<�0�<<��<{�<���<"K�<���<9��<D��<`   `   T�<��<wX�<?4�<���<�)�<���<�<��<Y��<���<�]�<V5�<�]�<���<Y��<��<�<���<�)�<���<?4�<wX�<��<`   `   ��<	A�<���<�m�<)�<�x�<Y��<he�<2�<��<�L�<��<ܯ�<��<�L�<��<2�<he�<Y��<�x�<)�<�m�<���<	A�<`   `   �r�<�6�<.��<{�<"&�<~��<�)�<O��<���<!��<���<_W�<�1�<_W�<���<!��<���<O��<�)�<~��<"&�<{�<.��<�6�<`   `   �B�<�
�<�i�<�n�<�1�<���<j�<�<���<��<vR�<���<��<���<vR�<��<���<�<j�<���<�1�<�n�<�i�<�
�<`   `   ��<��<JA�<�\�<�<�<W��<���<~��<�r�<���<Z��<���<�m�<���<Z��<���<�r�<~��<���<W��<�<�<�\�<JA�<��<`   `   ���<*��<$�<FX�<�W�<�8�<��<��<�
�<-B�<5��<IS�<65�<IS�<5��<-B�<�
�<��<��<�8�<�W�<FX�<$�<*��<`   `   Ƽ�<��<|"�<�p�<��<��<ݖ�<Z��<h��<��<ڍ�<�<�<� �<�<�<ڍ�<��<h��<Z��<ݖ�<��<��<�p�<|"�<��<`   `   ���<���<�I�<i��<���<~�<L<�<�f�<&��<�<��<zO�<�6�<zO�<��<�<&��<�f�<L<�<~�<���<i��<�I�<���<`   `   c�<���<��<� �<F�<��<��<�X�<9��<�/�<y��<R��<�y�<R��<y��<�/�<9��<�X�<��<��<F�<� �<��<���<`   `   '|�<ze�<�"�<B��<�6�<q��<?	�<v�<���<���<*2�<. �<���<. �<*2�<���<���<v�<?	�<q��<�6�<B��<�"�<ze�<`   `   ��<��<<��<H�<L�<���<�0�<��<J[�<��<���<���<���<���<���<��<J[�<��<�0�<���<L�<H�<<��<��<`   `   F��<&��<���<�i�<e!�<���<��<84�<���<%��<���<K}�<;v�<K}�<���<%��<���<84�<��<���<e!�<�i�<���<&��<`   `   v��<Ȫ�<Ô�<Lr�<yH�<��<���<���<��<מ�<C��<���<���<���<C��<מ�<��<���<���<��<xH�<Lr�<Ô�<Ȫ�<`   `   [��<��<̚�<Q��<*��<���<���<��<���<̫�<j��<:��<���<:��<j��<̫�<���<��<���<���<*��<Q��<̚�<��<`   `   %��<ץ�<��<ʽ�<4��<���<�*�<�c�<1��<���<'�<�&�<w2�<�&�<'�<���<1��<�c�<�*�<���<4��<ʽ�<��<ץ�<`   `   ��<έ�< ��<���<"-�<)}�<���<zE�<���<�<p�<O��<���<O��<p�<�<���<zE�<���<)}�<"-�<���< ��<έ�<`   `   R��<Q��<D��<��<@��<���<q��<
0�<��<j�<��<�1�<�L�<�1�<��<j�<��<
0�<q��<���<@��<��<C��<Q��<`   `   ە�<Ǩ�<���<�B�<���<�t�<�7�<U�<��<��<�K�<���<���<���<�K�<��<��<U�<�7�<�t�<���<�B�<���<Ǩ�<`   `   �x�<��<���<\T�<I��<���<��<���<���<���<���<��<�<�<��<���<���<���<���<��<���<H��<\T�<���<��<`   `   �F�<1d�<���<N�<��<��<:�<�u�<9��<���<ҩ�<�:�<�l�<�:�<ҩ�<���<9��<�u�<:�<��<��<N�<���<1d�<`   `   � �<�!�<R��<I,�<��<�.�<9|�<G��<0@�<{}�<�x�<��<?R�<��<�x�<{}�<0@�<G��<9|�<�.�<��<I,�<R��<�!�<`   `   ���<0��<�6�<��<��<� �<��<7�<���<���<���<"��<���<"��<���<���<���<7�<��<� �<��<��<�6�<0��<`   `   �6�<]�<���<���<���<"��<f�<O��<0��<e��<}�<���<��<���<}�<e��<0��<O��<f�<"��<���<���<���<]�<`   `   ߹�<��<�Y�<� �<�0�<<��<{�<���<"K�<���<9��<E��<C��<E��<9��<���<"K�<���<{�<<��<�0�<� �<�Y�<��<`   `   V5�<�]�<���<Z��<��<�<��<�)�<���<?4�<wX�<��<T�<��<wX�<?4�<���<�)�<���<�<��<Z��<���<�]�<`   `   ܯ�<��<�L�<��<2�<ie�<Y��<�x�<*�<�m�<���<	A�<��<	A�<���<�m�<*�<�x�<Y��<ie�<2�<��<�L�<��<`   `   �1�<_W�<���<!��<���<O��<�)�<~��<#&�<	{�</��<�6�<�r�<�6�</��<	{�<#&�<~��<�)�<O��<���<!��<���<_W�<`   `   ��<���<wR�<��<���<�<j�<���<�1�<�n�<�i�<�
�<�B�<�
�<�i�<�n�<�1�<���<j�<�<���<��<wR�<���<`   `   �m�<���<[��<���<�r�<��<���<X��<�<�<�\�<JA�<��<��<��<JA�<�\�<�<�<X��<���<��<�r�<���<[��<���<`   `   75�<JS�<5��<-B�<�
�<��<��<�8�<�W�<FX�<$�<+��<���<+��<$�<FX�<�W�<�8�<��<��<�
�<-B�<5��<JS�<`   `   K�<hm�<���<�x�<N]�<4p�<���<B�<VM�<�v�<�b�<{��<�.�<{��<�b�<�v�<VM�<A�<���<4p�<N]�<�x�<���<hm�<`   `   �f�<c��<���<Er�<�:�<�/�<y?�<�c�<��<���<�K�<7��<���<7��<�K�<���<��<�c�<y?�<�/�<�:�<Er�<���<c��<`   `   Թ�<���<�!�<��<�N�<� �<�<h��<���<w��<�p�<���<b�<���<�p�<w��<���<h��<�<� �<�N�<��<�!�<���<`   `   VJ�<``�<���<��<���<5K�<��<���<���<�H�<���<�,�<QK�<�,�<���<�H�<���<���<��<5K�<���<��<���<``�<`   `   I�<�/�<c�<_��<�$�<��<�D�<.��<��<S	�<Qv�<���<���<���<Qv�<S	�<��<.��<�D�<��<�$�<_��<c�<�/�<`   `   3�<
>�<}_�<���<���<D�<c��<��<���<J��<�D�<�x�<j��<�x�<�D�<J��<���<��<c��<D�<���<���<}_�<
>�<`   `   ���<[��<B��<��<��<��<9E�<���<O��<�<'8�<DZ�<rf�<DZ�<'8�<�<O��<���<9E�<��<��<��<B��<[��<`   `   �7�<�3�<�'�<��<��<Q��<���<-	�<��<�/�<�D�<9T�<�Y�<9T�<�D�<�/�<��<-	�<���<Q��<��<��<�'�<�3�<`   `   ��<M�<���<���<�\�<G�<���<��<m�<~i�<�^�<�Z�<�X�<�Z�<�^�<~i�<m�<��<���<G�<�\�<���<���<M�<`   `   ��<D��<3��<L�<x��<�B�<��<�F�<K��<է�<�z�<�b�<�Y�<�b�<�z�<է�<K��<�F�<��<�B�<x��<L�<3��<D��<`   `   �<���<���<^ �<�C�<�t�<��<���<�Q�<���<���<�a�<�R�<�a�<���<���<�Q�<���<��<�t�<�C�<^ �<���<���<`   `   ��<!��<m�<���<���<ؗ�<���<���<���<��<J��<$Q�<�:�<$Q�<J��<��<���<���<���<ؗ�<���<���<m�<!��<`   `   ��<P��<H�<�"�<w��<n��<kA�< �<M��<�<~��<I*�<G�<I*�<~��<�<M��< �<kA�<n��<w��<�"�<H�<P��<`   `   �u�<k6�<�}�<_�<K��<�e�<���<FS�<��<��<rU�<���<���<���<rU�<��<��<FS�<���<�e�<K��<_�<�}�<k6�<`   `   :��<�X�<ڈ�<SF�<���<���<u!�<�s�<���<���<��<_��<�a�<_��<��<���<���<�s�<u!�<���<���<SF�<ڈ�<�X�<`   `   ZW�<8	�<(�<4��<��<a%�<�1�<\�<5��<}�<ԕ�<��<���<��<ԕ�<}�<5��<\�<�1�<a%�<��<4��<(�<8	�<`   `   ��<A�<JT�<���<�<�
�<��<}
�<�Z�<k�<�	�<�}�<�L�<�}�<�	�<k�<�Z�<}
�<��<�
�<�<���<JT�<A�<`   `   yS�<���<��<J��<u��<ޠ�<t��<��<���<�g�<�i�<��<,��<��<�i�<�g�<���<��<t��<ޠ�<u��<J��<��<���<`   `   ���<O�<*[�<<��<&�<T��<]��<���<&�<��<*��<1(�<���<1(�<*��<��<&�<���<]��<T��<&�<<��<*[�<O�<`   `   ���<�?�<�Q�<���<��<��<���<��<vX�<���<��<�x�<bG�<�x�<��<���<vX�<��<���<��<��<���<�Q�<�?�<`   `   8�<��<(�<d��<���<��<��<,-�<v��<�G�<�a�<"��<?��<"��<�a�<�G�<v��<,-�<��<��<���<d��<(�<��<`   `   e��<kj�<���<�M�<ů�<���<:�<�T�<��<՟�<���<�C�<�<�C�<���<՟�<��<�T�<:�<���<ů�<�M�<���<kj�<`   `   ��<���<��<<��<�s�<���<`!�<:��<g.�<H�<�M�<���<6��<���<�M�<H�<g.�<:��<_!�<���<�s�<<��<��<���<`   `   l��<6Y�<	��<���<�L�<	��<S�<���<5��<k��<K��<���<�c�<���<K��<k��<5��<���<S�<	��<�L�<���<	��<6Y�<`   `   �.�<{��<�b�<�v�<VM�<A�<���<4p�<M]�<�x�<���<hm�<K�<hm�<���<�x�<M]�<4p�<���<A�<VM�<�v�<�b�<{��<`   `   ���<6��<�K�<���<��<�c�<y?�<�/�<�:�<Er�<���<b��<�f�<b��<���<Er�<�:�<�/�<y?�<�c�<��<���<�K�<6��<`   `   a�<���<�p�<w��<���<g��<�<� �<�N�<��<�!�<���<ӹ�<���<�!�<��<�N�<� �<�<g��<���<w��<�p�<���<`   `   PK�<�,�<���<�H�<���<���<��<5K�<���<��<���<_`�<UJ�<_`�<���<��<���<5K�<��<���<���<�H�<���<�,�<`   `   ���<���<Qv�<S	�<��<.��<�D�<��<�$�<_��<c�<�/�<H�<�/�<c�<_��<�$�<��<�D�<.��<��<S	�<Qv�<���<`   `   j��<�x�<�D�<J��<���<��<c��<D�<���<���<}_�<	>�<3�<	>�<}_�<���<���<D�<c��<��<���<J��<�D�<�x�<`   `   rf�<DZ�<'8�<�<O��<���<9E�<��<��<��<B��<Z��<���<Z��<B��<��<��<��<9E�<���<O��<�<'8�<DZ�<`   `   �Y�<9T�<�D�<�/�<��<,	�<���<Q��<��<��<�'�<�3�<�7�<�3�<�'�<��<��<Q��<���<,	�<��<�/�<�D�<9T�<`   `   �X�<�Z�<�^�<~i�<m�<��<���<G�<�\�<���<���<M�<��<M�<���<���<�\�<G�<���<��<m�<~i�<�^�<�Z�<`   `   �Y�<�b�<�z�<է�<J��<�F�<��<�B�<x��<L�<3��<C��<��<C��<3��<L�<x��<�B�<��<�F�<J��<է�<�z�<�b�<`   `   �R�<�a�<���<���<�Q�<���<��<�t�<�C�<^ �<���<���<�<���<���<^ �<�C�<�t�<��<���<�Q�<���<���<�a�<`   `   �:�<$Q�<J��<��<���<���<���<ؗ�<���<���<m�<!��<��<!��<m�<���<���<ؗ�<���<���<���<��<J��<$Q�<`   `   G�<I*�<~��<�<M��< �<kA�<n��<w��<�"�<H�<P��<��<P��<H�<�"�<w��<n��<jA�< �<M��<�<~��<I*�<`   `   ���<���<rU�<��<��<GS�<���<�e�<K��<_�<�}�<k6�<�u�<k6�<�}�<_�<K��<�e�<���<FS�<��<��<rU�<���<`   `   �a�<_��<��<���<���<�s�<u!�<���<���<SF�<ڈ�<�X�<:��<�X�<ڈ�<SF�<���<���<u!�<�s�<���<���<��<_��<`   `   ���<��<ԕ�<}�<5��<\�<�1�<b%�<��<4��<(�<8	�<ZW�<8	�<(�<4��<��<b%�<�1�<\�<5��<}�<ԕ�<��<`   `   �L�<�}�<�	�<k�<�Z�<}
�<��<�
�<�<���<KT�<A�<��<A�<KT�<���<�<�
�<��<}
�<�Z�<k�<�	�<�}�<`   `   ,��< ��<�i�<�g�<���<��<t��<ޠ�<v��<K��<��<���<yS�<���<��<K��<v��<ޠ�<t��<��<���<�g�<�i�< ��<`   `   ���<1(�<*��<��<'�<���<^��<U��<'�<<��<*[�<O�<���<O�<*[�<<��<'�<U��<^��<���<&�<��<*��<1(�<`   `   cG�<�x�<��<���<vX�<��<���<��<��<���<�Q�<�?�<���<�?�<�Q�<���<��<��<���<��<vX�<���<��<�x�<`   `   ?��<"��<�a�<�G�<v��<,-�<��<��<���<e��<(�<��<8�<��<(�<e��<���<��<��<,-�<v��<�G�<�a�<"��<`   `   �<�C�<���<֟�<��<�T�<:�<���<ů�<�M�<���<kj�<f��<kj�<���<�M�<ů�<���<:�<�T�<��<֟�<���<�C�<`   `   6��<���<�M�<I�<h.�<;��<`!�<���<�s�<<��<��<���<��<���<��<<��<�s�<���<`!�<;��<h.�<I�<�M�<���<`   `   �c�<���<L��<l��<5��<���<S�<	��<�L�<���<	��<6Y�<l��<6Y�<	��<���<�L�<	��<S�<���<5��<l��<L��<���<`   `   p��<��<l��<Y�<t�<���<hb�<Z	�<���<��<�=�<��<i:�<��<�=�<��<���<Z	�<gb�<���<t�<Y�<l��<��<`   `   ��<4�<���<`[�<2Q�<Ǉ�<���<�Z�<���<�<Y�<O��<���<O��<Y�<�<���<�Z�<���<Ǉ�<2Q�<`[�<���<4�<`   `   �s�<ޔ�<g��<���<hx�<N��<L��<���<�$�<G9�<)�</��<���</��<)�<G9�<�$�<���<L��<N��<hx�<���<f��<ޔ�<`   `   s�<0:�<���</�<���<"��<���<��<���<A��<�f�<���<T�<���<�f�<A��<���<��<���<"��<���</�<���<0:�<`   `   P�<6�<�{�<���<_��<�=�<��<��<L��<�j�<f��<|[�<�{�<|[�<f��<�j�<L��<��<��<�=�<^��<���<�{�<6�<`   `   v�<'��<��<N
�<dx�<e��<!��<o:�<���<�_�<$��<_�<�-�<_�<$��<�_�<���<o:�<!��<e��<dx�<N
�<��<'��<`   `   �"�<�+�<�D�<�p�<C��<T��<�T�<���<+#�<��<,��<���<&�<���<,��<��<+#�<���<�T�<T��<C��<�p�<�D�<�+�<`   `   �<��<��<��<h�<*�<'@�<S`�<���<q��<���<T �<�	�<T �<���<q��<���<S`�<'@�<*�<h�<��<��<��<`   `   R�<�F�<Z&�<��<���<'��<�J�<Y"�<�	�<���<��<`
�<��<`
�<��<���<�	�<Y"�<�J�<'��<���<��<Z&�<�F�<`   `   ۰�<E��<hW�<K��<�s�<���<Ed�<���<��<OK�<�%�<��<�
�<��<�%�<OK�<��<���<Ed�<���<�s�<K��<hW�<E��<`   `   ��<���<+��<k��<=/�<6V�<I|�<���<��<ڋ�<~4�<v	�<���<v	�<~4�<ڋ�<��<���<I|�<6V�<=/�<k��<+��<���<`   `   �z�<J�<���<V��<���<��<Q}�<�d�<�r�<���<�1�<���<G��<���<�1�<���<�r�<�d�<Q}�<��<���<V��<���<J�<`   `   I��<�d�< ��<l��<�M�<#��<=S�<��<���<���<��<��<S��<��<��<���<���<��<=S�<#��<�M�<l��< ��<�d�<`   `   p�<�(�<"Y�<p�<0}�<η�<��<�@�<%��<��< ��<�F�<�#�<�F�< ��<��<%��<�@�<��<η�<0}�<p�<"Y�<�(�<`   `   ���<+{�<0��<A�<�O�<�J�<y?�<�T�<���<�M�<�T�<���<e��<���<�T�<�M�<���<�T�<y?�<�J�<�O�<A�<0��<+{�<`   `   ؠ�<H�<F�<4��<���<�~�<??�<�#�<�K�<���<���<��<N��<��<���<���<�K�<�#�<??�<�~�<���<4��<F�<H�<`   `   c��<���<�u�<d��<���<�P�<7��<&��<��<�#�<���<\P�<�<\P�<���<�#�<��<&��<7��<�P�<���<d��<�u�<���<`   `   ؜�<�:�<��<d�<�5�<X��<0O�<���<���<�U�<�&�<Sr�<N<�<Sr�<�&�<�U�<���<���<0O�<X��<�5�<d�<��<�:�<`   `   &��<Cn�<�O�<��<�^�<C��<	q�<��<�<�n�<?�<��<FT�<��<?�<�n�<�<��<	q�<C��<�^�<��<�O�<Cn�<`   `   p��<^6�<V�<Ce�<Y;�<��<�e�<��<+�<�~�<�U�<��<�p�<��<�U�<�~�<+�<��<�e�<��<Y;�<Ce�<V�<^6�<`   `   6�<I��<|��<���<%��<���<�A�<t�<�"�<���<�y�<���<[��<���<�y�<���<�"�<t�<�A�<���<%��<���<|��<I��<`   `   �P�<��<���<�k�<By�<fO�<��<��<Z9�<���<t��<@ �<���<@ �<t��<���<Z9�<��<��<fO�<By�<�k�<���<��<`   `   +��<,4�<�H�<P��<��</�<	�<��<�p�<�<]!�<���<�c�<���<\!�<�<�p�<��<	�</�<��<P��<�H�<,4�<`   `   p��<���<���<�d�<���<���<�<�\�<>��<��<r��<t9�<��<t9�<r��<��<>��<�\�<�<���<���<�d�<���<���<`   `   h:�<��<�=�<��<���<Z	�<gb�<���<t�<Y�<k��<��<o��<��<k��<Y�<t�<���<gb�<Z	�<���<��<�=�<��<`   `   ���<N��<X�<�<���<�Z�<���<Ǉ�<2Q�<`[�<���<4�<��<4�<���<`[�<2Q�<Ƈ�<���<�Z�<���<�<X�<N��<`   `   ���<.��<(�<G9�<�$�<���<K��<M��<hx�<���<f��<ޔ�<�s�<ݔ�<f��<���<hx�<M��<K��<���<�$�<G9�<(�<.��<`   `   S�<���<�f�<@��<���<��<���<!��<���</�<���<0:�<s�<0:�<���</�<���<!��<���<��<���<@��<�f�<���<`   `   �{�<|[�<f��<�j�<L��<��<��<�=�<^��<���<�{�<6�<O�<6�<�{�<���<^��<�=�<��<��<L��<�j�<f��<|[�<`   `   �-�<^�<$��<�_�<���<o:�<!��<e��<dx�<M
�<��<&��<v�<&��<��<M
�<dx�<e��<!��<o:�<���<�_�<$��<^�<`   `   %�<���<+��<��<+#�<���<�T�<S��<B��<�p�<�D�<�+�<�"�<�+�<�D�<�p�<B��<S��<�T�<���<+#�<��<+��<���<`   `   �	�<T �<���<q��<���<S`�<'@�<*�<g�<��<��<��<�<��<��<��<g�<*�<&@�<S`�<���<p��<���<T �<`   `   ��<`
�<��<���<�	�<Y"�<�J�<'��<���<��<Z&�<�F�<R�<�F�<Z&�<��<���<'��<�J�<X"�<�	�<���<��<`
�<`   `   �
�<��<�%�<NK�<��<���<Ed�<���<�s�<J��<hW�<E��<ڰ�<E��<hW�<J��<�s�<���<Ed�<���<��<NK�<�%�<��<`   `   ���<v	�<~4�<ڋ�<��<���<I|�<6V�<=/�<k��<+��<���<��<���<+��<k��<=/�<6V�<I|�<���<��<ڋ�<~4�<u	�<`   `   G��<���<�1�<���<�r�<�d�<Q}�<��<���<V��<���<J�<�z�<J�<���<V��<���<��<Q}�<�d�<�r�<���<�1�<���<`   `   S��<��<��<���<���<��<=S�<#��<�M�<l��< ��<�d�<I��<�d�<��<l��<�M�<#��<=S�<��<���<���<��<��<`   `   �#�<�F�<��<��<%��<�@�<��<η�<0}�<p�<"Y�<�(�<p�<�(�<"Y�<p�<0}�<η�<��<�@�<$��<��< ��<�F�<`   `   e��<���<�T�<�M�<���<�T�<y?�<�J�<�O�<A�<1��<+{�<���<+{�<0��<A�<�O�<�J�<y?�<�T�<���<�M�<�T�<���<`   `   N��<��<���<���<�K�<�#�<??�<�~�<���<5��<F�<H�<ؠ�<H�<F�<5��<���<�~�<??�<�#�<�K�<���<���<��<`   `   �<\P�<���<�#�<��<&��<7��< Q�<���<e��<�u�<���<c��<���<�u�<d��<���<�P�<7��<&��<��<�#�<���<\P�<`   `   N<�<Tr�<�&�<�U�<���<���<1O�<X��<�5�<d�<��<�:�<؜�<�:�<��<d�<�5�<X��<1O�<���<���<�U�<�&�<Tr�<`   `   GT�<��<?�<�n�<�<��<	q�<D��<�^�<��<�O�<Cn�<'��<Cn�<�O�<��<�^�<D��<	q�<��<�<�n�<?�<��<`   `   �p�<��<�U�<�~�<,�<��<�e�<��<Z;�<Ce�<W�<_6�<p��<_6�<W�<Ce�<Z;�<��<�e�<��<,�<�~�<�U�<��<`   `   [��<���<�y�<���<�"�<t�<�A�<���<%��<���<}��<I��<7�<I��<}��<���<%��<���<�A�<t�<�"�<���<�y�<���<`   `   ���<A �<u��<���<Z9�<��<��<gO�<By�<�k�<���<��<�P�<��<���<�k�<By�<gO�<��<��<Z9�<���<u��<A �<`   `   �c�<���<]!�<�<�p�<��<	�</�<��<Q��<�H�<,4�<+��<,4�<�H�<Q��<��</�<	�<��<�p�<�<]!�<���<`   `   ��<t9�<s��<��<?��<�\�<�<���<���<�d�<���< ��<q��< ��<���<�d�<���<���<�<�\�<?��<��<s��<t9�<`   `   
��<��<?��<���<���<n�<2�<��<��<�v�<���<��<���<��<���<�v�<��<��<2�<n�<���<���<?��<��<`   `   �<�B�<G��<��<(��<qB�<~��<l��<�0�<���<���<��<i��<��<���<���<�0�<l��<~��<pB�<(��<��<G��<�B�<`   `   ��<N��<�*�<B��<+	�<�]�<���<�S�<���<��<'�<���<���<���<&�<��<���<�S�<���<�]�<+	�<B��<�*�<N��<`   `   �E�<Gm�<s��<e��<���<ٹ�<\�<�Y�<���<��<���<H$�<!U�<H$�<���<��<���<�Y�<\�<ٹ�<���<e��<s��<Gm�<`   `   �_�<���<���<���<�d�<_�<�w�<1��<I��<O��<	U�<���<^��<���<	U�<O��<I��<1��<�w�<_�<�d�<���<���<���<`   `   ���<,��<�>�<S��<�w�<�H�<�&�<��<u��<b��<�B�<ѣ�<���<ѣ�<�B�<b��<t��<��<�&�<�H�<�w�<S��<�>�<,��<`   `   ]��<��<���<|E�<j��<c�<
�<���<�O�<���<�T�<R��<���<R��<�T�<���<�O�<���<
�<c�<j��<|E�<���<��<`   `   ��<ם�<���<��<^L�<Ǩ�<��<�s�<���<#1�<*{�<���<��<���<*{�<#1�<���<�s�<��<Ǩ�<^L�<��<���<ם�<`   `   T��<���<���<���<?��<��<�%�<�D�<�d�<Y��<���<P��<���<P��<���<Y��<�d�<�D�<�%�<��<?��<���<���<���<`   `   �6�<',�<��<���<6��<�x�<�B�<��<y��<��<B��<k��<���<k��<B��<��<y��<��<�B�<�x�<6��<���<��<',�<`   `   ���<���<�K�<t��<'i�<���<�Q�<���<�a�<�
�<]��<y��<T��<y��<]��<�
�<�a�<���<�Q�<���<'i�<t��<�K�<���<`   `   ���<)��<�o�<���<w�<�#�<�?�<@j�<J��<��<���<Ms�<�X�<Ms�<���<��<J��<@j�<�?�<�#�<w�<���<�o�<)��<`   `   ��<���<`[�<~�<�f�<n2�<��<���<V��<$�<$l�<a�<���<a�<$l�<$�<U��<���<��<n2�<�f�<~�<`[�<���<`   `   ���<~��<N��<���<|�<���<n�<1��<Ƿ�<?��<`��<���<bT�<���<`��<?��<Ƿ�<1��<n�<���<|�<���<N��<~��<`   `   {"�<��<��<���<k0�<$c�<��<���<K]�<�)�<VH�<"��<���<"��<VH�<�)�<K]�<���<��<$c�<k0�<���<��<��<`   `   ���<���<v��<G�<�w�<o�<�`�<s�<l��<j�<�l�<C��<��<C��<�l�<j�<l��<s�<�`�<o�<�w�<G�<u��<���<`   `   �'�<���<[��<'H�<P�<x�<o��<`��<0��<z�<�h�<P��<���<P��<�h�<z�<0��<`��<o��<x�<P�<'H�<[��<���<`   `   a��<	��<e{�<���<���<�m�<�<���<F��<6g�<1H�< ��<~[�< ��<1H�<6g�<F��<���<�<�m�<���<���<e{�<	��<`   `   �*�<��<��<<�<���<�y�<��<���<u��<0B�<�<5k�< +�<5k�<�<0B�<u��<���<��<�y�<���<<�<��<��<`   `   W�<g��<
��<���<���<�U�<���<'��<���<u�<+��<:D�<��<:D�<+��<u�<���<'��<���<�U�<���<���<
��<g��<`   `   ���<T�<�>�<\��<'q�<��<���<��<Д�<��<���<�7�<���<�7�<���<��<Д�<��<���<��<'q�<\��<�>�<T�<`   `   �+�<���<��<�&�<��<N��<3��<�t�<d��<�<a��<�V�<N�<�V�<a��<�<d��<�t�<3��<N��<��<�&�<��<���<`   `   ���<nE�<YJ�<���<��<L��<��<)��<���<UW�<�K�<Y��<�|�<Y��<�K�<UW�<���<)��<��<L��<��<���<YJ�<nE�<`   `   �$�<*��<���<��<]��<Y��<���<���<o1�<F��<r��<�?�<��<�?�<r��<F��<o1�<���<���<Y��<]��<��<���<*��<`   `   ���<��<���<�v�<��<��<2�<n�<���<���<?��<��<
��<��<?��<���<���<n�<2�<��<��<�v�<���<��<`   `   i��<��<���<���<�0�<k��<~��<pB�<(��<��<F��<�B�<�<�B�<F��<��<(��<pB�<~��<k��<�0�<���<���<��<`   `   ���<���<&�<��<���<�S�<���<�]�<+	�<A��<�*�<N��<��<N��<�*�<A��<+	�<�]�<���<�S�<���<��<&�<���<`   `    U�<H$�<���<��<���<�Y�<[�<ع�<���<e��<s��<Gm�<�E�<Gm�<s��<e��<���<ع�<[�<�Y�<���<��<���<H$�<`   `   ]��<���<U�<N��<H��<0��<�w�<_�<�d�<���<���<���<�_�<���<���<���<�d�<_�<�w�<0��<H��<N��<U�<���<`   `   ���<У�<�B�<a��<t��<��<�&�<�H�<�w�<S��<�>�<+��<���<+��<�>�<S��<�w�<�H�<�&�<��<t��<a��<�B�<У�<`   `   ���<R��<�T�<���<�O�<���<
�<c�<j��<|E�<���<��<\��<��<���<|E�<j��<c�<
�<���<�O�<���<�T�<R��<`   `   ��<���<){�<#1�<���<�s�<��<Ǩ�<^L�<��<���<֝�<��<֝�<���<��<^L�<Ǩ�<��<�s�<���<#1�<){�<���<`   `   ���<P��<���<X��<�d�<�D�<�%�<��<?��<���<���<���<S��<���<���<���<>��<��<�%�<�D�<�d�<X��<���<P��<`   `   ���<k��<B��<��<y��<��<�B�<�x�<6��<���<��<&,�<�6�<&,�<��<���<5��<�x�<�B�<��<y��<��<A��<k��<`   `   T��<y��<]��<�
�<�a�<���<�Q�<���<'i�<t��<�K�<���<���<���<�K�<t��<&i�<���<�Q�<���<�a�<�
�<]��<y��<`   `   �X�<Ms�<���<��<J��<@j�<�?�<�#�<w�<���<�o�<)��<���<)��<�o�<���<w�<�#�<�?�<@j�<J��<��<���<Ms�<`   `   ���<a�<$l�<$�<V��<���<��<n2�<�f�<~�<`[�<���<��<���<`[�<~�<�f�<n2�<��<���<U��<$�<$l�<a�<`   `   bT�<���<`��<?��<Ƿ�<1��<n�<���<|�<���<N��<~��<���<~��<N��<���<|�<���<n�<1��<Ƿ�<?��<`��<���<`   `   ���<"��<VH�<�)�<K]�<���<��<$c�<k0�<���<��<��<{"�<��<��<���<k0�<$c�<��<���<K]�<�)�<VH�<"��<`   `   ��<C��<�l�<j�<l��<s�<�`�<o�<�w�<G�<v��<���<���<���<v��<G�<�w�<o�<�`�<s�<l��<j�<�l�<C��<`   `   ���<P��<�h�<z�<0��<`��<o��<x�<P�<(H�<[��<���<�'�<���<[��<(H�<P�<x�<o��<`��<0��<z�<�h�<P��<`   `   ~[�< ��<1H�<7g�<G��<���<�<�m�<���<���<e{�<	��<b��<	��<e{�<���<���<�m�<�<���<F��<7g�<1H�< ��<`   `    +�<6k�<�<1B�<v��<���<��<�y�<���<<�<��<��<�*�<��<��<<�<���<�y�<��<���<v��<1B�<�<6k�<`   `   ��<:D�<,��<v�<���<'��<���<�U�<���< ��<��<h��<W�<h��<��< ��<���<�U�<���<'��<���<v�<,��<:D�<`   `   ���<�7�<���<��<Д�<��<���<��<(q�<]��<�>�<T�<���<T�<�>�<]��<'q�<��<���<��<Д�<��<���<�7�<`   `   O�<�V�<b��<�<d��<�t�<4��<O��<��<�&�<��<���<�+�<���<��<�&�<��<O��<3��<�t�<d��<�<b��<�V�<`   `   �|�<Y��<�K�<UW�<���<)��<��<M��<��<���<ZJ�<oE�<���<oE�<ZJ�<���<��<M��<��<)��<���<UW�<�K�<Y��<`   `   ��<�?�<s��<G��<p1�<���<���<Z��<^��<��<���<+��<�$�<+��<���<��<^��<Y��<���<���<o1�<G��<s��<�?�<`   `   a(�<a^�<���<6��<�<m��<�+�<���<�~�<)��<��<)��<��<)��<��<)��<�~�<���<�+�<m��<�<6��<���<a^�<`   `   yX�<��<��<3�<NY�<���< z�<�"�<���<��<"7�<���<�&�<���<"7�<��<���<�"�< z�<���<NY�<3�<��<��<`   `   a��<���<���<֑�<K��<~[�<f��<[��<
�<�l�<(s�<��<�S�<��<(s�<�l�<	�<[��<e��<~[�<K��<֑�<���<���<`   `   Sj�<���<�?�<B�<`��<U�<���<�(�<���<H��<+��<`�<ߔ�<`�<+��<G��<���<�(�<���<U�<`��<B�<�?�<���<`   `   MJ�<��<}#�<l�<�d�<���<�[�<d��<�&�<sE�<|%�<��<���<��<|%�<rE�<�&�<d��<�[�<���<�d�<l�<}#�<��<`   `   ]�<��<�-�<#�<�V�<���<�%�<��<���<r��< ��<O��<3(�<O��< ��<r��<���<��<�%�<���<�V�<#�<�-�<��<`   `   5��<C��<*`�<�D�<]f�<��<���<�1�<�H�<�-�<E��<�>�<Xh�<�>�<E��<�-�<�H�<�1�<���<��<]f�<�D�<*`�<C��<`   `   � �<g.�<n��<��<5��<!��<���<���<���<&��<��<jr�<��<jr�<��<&��<���<���<���<!��<5��<��<n��<g.�<`   `   -�<��<��<Y��<���<��<b��<#q�<S:�<��<�H�<���<���<���<�H�<��<S:�<#q�<b��<��<���<Y��<��<��<`   `   -��<��<H~�<)�<���<i{�<:�<2��<a��<� �<IX�<*��<��<*��<IX�<� �<a��<2��<:�<i{�<���<)�<H~�<��<`   `   �b�<�}�<M��<�8�<ۼ�<�C�<���<�?�<[��<���<�4�<SP�<�Z�<SP�<�4�<���<[��<�?�<���<�C�<ۼ�<�8�<M��<�}�<`   `   '��<��<���<�2�<���<\��<�"�<�^�<6��<���<^��<���<<��<���<^��<���<6��<�^�<�"�<\��<���<�2�<���<��<`   `   ���<���<���< ��<j�<%6�<�A�<dA�<�A�<B�<D�<�A�<UB�<�A�<D�<B�<�A�<dA�<�A�<%6�<j�< ��<���<���<`   `   E1�<9�<�L�<�^�<	_�<<H�<h�<���<���<��<�o�<�_�<�[�<�_�<�o�<��<���<���<h�<<H�<	_�<�^�<�L�<9�<`   `   [��<���<��<ш�<N^�<��<��<�A�<��<��<I]�<6C�<|<�<6C�<I]�<��<��<�A�<��<��<N^�<ш�<��<���<`   `   /��<:��<n��<�u�<+�<��<��<�d�<��<Md�<��<���<U��<���<��<Md�<��<�d�<��<��<+�<�u�<n��<:��<`   `   ���<W��<v��<�4�<���<<��<,�<�Y�<���<��<���<-�<q�<-�<���<��<���<�Y�<,�<<��<���<�4�<v��<W��<`   `   G��<9��<Z�<���<�<;5�<b3�<�3�<�S�<~��<2�<���<��<���<2�<~��<�S�<�3�<b3�<;5�<�<���<Z�<9��<`   `   '��<���<��<m�<^��<dd�<2�<��<��<�@�<A��<bn�<�X�<bn�<A��<�@�<��<��<2�<cd�<^��<m�<��<���<`   `   І�<&Z�<���<a�<���<V��<};�<���<��<���<bX�<@��<���<@��<bX�<���<��<���<};�<V��<���<a�<���<&Z�<`   `   Lh�<�2�<���<��<gY�<���<Ac�<x��<��<���<<!�<��<���<��<<!�<���<��<x��<Ac�<���<gY�<��<���<�2�<`   `   5I�<V�<4^�<�I�<���<nV�<'��</6�<,��<-��<!&�<ű�<���<ű�<!&�<-��<,��</6�<'��<nV�<���<�I�<4^�<V�<`   `   -�<:��< 3�<O�<���<h��<EH�<���<8Y�<+?�<�r�<T��<r��<T��<�r�<+?�<8Y�<���<EH�<h��<���<O�< 3�<:��<`   `   e�<���<��<m��<�t�<~��<��<�}�<8�<8��<(�<׆�<�S�<׆�<(�<8��<8�<�}�<��<~��<�t�<m��<��<���<`   `   ��<(��<��<(��<�~�<���<�+�<l��<�<6��<���<a^�<`(�<`^�<���<6��<�<l��<�+�<���<�~�<(��<��<(��<`   `   �&�<���<!7�<��<���<�"�<�y�<���<NY�<3�<��<��<xX�<��<��<2�<NY�<���<�y�<�"�<���<��<!7�<���<`   `   �S�<��<'s�<�l�<	�<Z��<e��<}[�<J��<Ց�<���<���<`��<���<���<Ց�<J��<}[�<e��<Z��<	�<�l�<'s�<��<`   `   ޔ�<`�<*��<G��<���<�(�<���<T�<_��<B�<�?�<���<Rj�<���<�?�<B�<_��<T�<���<�(�<���<G��<*��<`�<`   `   ���<��<|%�<rE�<�&�<d��<�[�<���<�d�<l�<|#�<��<MJ�<��<|#�<l�<�d�<���<�[�<d��<�&�<rE�<|%�<��<`   `   2(�<O��< ��<q��<���<��<�%�<���<�V�< #�<�-�<��<]�<��<�-�< #�<�V�<���<�%�<��<���<q��< ��<O��<`   `   Wh�<�>�<D��<�-�<�H�<�1�<���<��<\f�<�D�<*`�<B��<5��<B��<*`�<�D�<\f�<��<���<�1�<�H�<�-�<D��<�>�<`   `   ��<jr�<��<%��<���<���<���< ��<5��<��<m��<g.�<� �<g.�<m��<��<5��< ��<���<���<���<%��<��<jr�<`   `   ���<���<�H�<��<S:�<"q�<a��<��<���<Y��<��<��<,�<��<��<Y��<���<��<a��<"q�<S:�<��<�H�<���<`   `   ��<)��<IX�<� �<a��<2��<
:�<i{�<���<)�<G~�<��<-��<��<G~�<)�<���<i{�<
:�<2��<a��<� �<IX�<)��<`   `   �Z�<RP�<�4�<���<[��<�?�<���<�C�<ۼ�<�8�<M��<�}�<�b�<�}�<M��<�8�<ۼ�<�C�<���<�?�<Z��<���<�4�<RP�<`   `   <��<���<^��<���<6��<�^�<�"�<\��<���<�2�<���<��<'��<��<���<�2�<���<\��<�"�<�^�<5��<���<^��<���<`   `   UB�<�A�<D�<B�<�A�<dA�<�A�<%6�<k�< ��<���<���<���<���<���< ��<j�<$6�<�A�<dA�<�A�<B�<D�<�A�<`   `   �[�<�_�<�o�<��<���<���<i�<<H�<
_�<�^�<�L�<9�<E1�<9�<�L�<�^�<	_�<<H�<h�<���<���<��<�o�<�_�<`   `   |<�<6C�<I]�<��<��<�A�<��<��<N^�<҈�<��<���<[��<���<��<ш�<N^�<��<��<�A�<��<��<I]�<6C�<`   `   V��<���<��<Nd�<��<�d�<��<��<+�<�u�<o��<:��</��<:��<n��<�u�<+�<��<��<�d�<��<Md�<��<���<`   `   q�<-�<���<��<���<�Y�<,�<<��<���<�4�<w��<W��<���<W��<v��<�4�<���<<��<,�<�Y�<���<��<���<-�<`   `   ��<���<2�<��<�S�<�3�<b3�<;5�<�<���<Z�<9��<G��<9��<Z�<���<�<;5�<b3�<�3�<�S�<~��<2�<���<`   `   �X�<cn�<B��<�@�<��<��<2�<dd�<_��<m�<��<���<(��<���<��<m�<^��<dd�<2�<��<��<�@�<A��<cn�<`   `   ���<@��<cX�<���<��<���<~;�<V��<���<b�<���<'Z�<ц�<'Z�<���<b�<���<V��<};�<���<��<���<cX�<@��<`   `   ���<��<<!�<���<��<x��<Bc�<���<hY�<��<���<�2�<Lh�<�2�<���<��<gY�<���<Ac�<x��<��<���<<!�<��<`   `   ���<ű�<!&�<-��<-��<06�<(��<oV�<���<�I�<5^�<W�<6I�<W�<5^�<�I�<���<nV�<(��<06�<-��<-��<!&�<ű�<`   `   s��<U��<�r�<,?�<8Y�<���<FH�<i��<���<P�<3�<;��<-�<;��< 3�<O�<���<i��<EH�<���<8Y�<,?�<�r�<U��<`   `   �S�<؆�<)�<9��<9�<�}�<��<~��<�t�<n��<��<���<f�<���<��<n��<�t�<~��<��<�}�<9�<9��<(�<؆�<`   `   '��<=��<X�<u��<�:�<���<���<C�<w%�<���<}�<�C�<�V�<�C�<}�<���<w%�<B�<���<���<�:�<u��<X�<=��<`   `   ��<D��<#l�<�@�<G�<"f�<���<à�<��<�l�<��<de�<Յ�<de�<��<�l�<��<à�<���<"f�<G�<�@�<"l�<D��<`   `   ���<R�<\��<���<�P�<��<dJ�<9��<��<O��<J��<V�<ZD�<V�<I��<O��<��<8��<dJ�<��<�P�<���<\��<Q�<`   `   ���<6:�<�#�<7��<N4�<��<���<�}�<���<D�<���<�j�<V��<�j�<���<D�<���<�}�<���<��<N4�<7��<�#�<6:�<`   `   ���<F�<sK�<��<���<Q��<'�<���<ؖ�<Y��<���<�Q�<@�<�Q�<���<Y��<ז�<���<'�<P��<���<��<sK�<F�<`   `   ���<�!�<A�<��<�0�<Ѝ�<���<�<m��<�9�<N4�<���<���<���<M4�<�9�<m��<�<���<Ѝ�<�0�<��<A�<�!�<`   `   #X�<���<���<���<|6�<��<�Q�<��<��<>!�<m0�<m��<���<m��<m0�<>!�<��<��<�Q�<��<|6�<���<���<���<`   `   ��<��<Ml�<�q�<Q��<��<�Z�<#��<P��<s��<w��<�c�<.��<�c�<w��<s��<P��<#��<�Z�<��<Q��<�q�<Ml�<��<`   `   ��<��<Nz�<���<yS�<D6�<�<���<���<��<[��<��<���<��<[��<��<���<���<�<D6�<yS�<���<Nz�<��<`   `   ���<1��<��<�s�<�U�<�i�<�i�<#�<�u�< G�<���<:a�<I��<:a�<���< G�<�u�<#�<�i�<�i�<�U�<�s�<��<1��<`   `   ;��<kw�<�2�<N��<��<9A�<Wp�<:K�<���<<��<��<���<�.�<���<��<<��<���<:K�<Wp�<9A�<��<N��<�2�<kw�<`   `   _Y�<n�<p��<��<�.�<n��<�#�<O$�<K��<��<G!�<?�<�_�<?�<G!�<��<K��<O$�<�#�<n��<�.�<��<p��<n�<`   `   ��<�V�<sg�<�{�<�&�<��<4��<-��<]N�<�b�<[��<���<`=�<���<[��<�b�<]N�<-��<4��<��<�&�<�{�<sg�<�V�<`   `   N��<=��<���<"(�<��<	�<��<K�<��<���<�l�<@s�<��<@s�<�l�<���<��<K�<��<	�<��<"(�<���<=��<`   `   ֠�<�m�<���<��<X�<m!�<?��<�>�<���<��<���<��<��<��<���<��<���<�>�<?��<m!�<X�<��<���<�m�<`   `   �<C��<6�<�r�<�e�<zs�<�7�<Qu�<u�<�0�<^��<A��<82�<A��<^��<�0�<u�<Qu�<�7�<zs�<�e�<�r�<6�<C��<`   `   w�<�9�<�`�<���<�T�<�-�<l��<���<�N�<J�<p��<���<8-�<���<p��<J�<�N�<���<l��<�-�<�T�<���<�`�<�9�<`   `   ��<���<G��<{��<���<�r�<���<�k�<���<dx�<���< ��<S$�< ��<���<dx�<���<�k�<���<�r�<���<{��<G��<���<`   `   f��<�Q�<,��<bz�<�a�<-W�<,�<Re�<uN�<��<;�<���<�1�<���<;�<��<uN�<Re�<,�<-W�<�a�<bz�<,��<�Q�<`   `   �n�<&��<@@�<�9�<���<���<��<���<{K�<h��<T��<�5�<_s�<�5�<T��<h��<{K�<���<��<���<���<�9�<@@�<&��<`   `   1��<5>�<8�<���<�H�<^��<�f�<��<t��<���<,J�<g��<���<g��<,J�<���<t��<��<�f�<^��<�H�<���<8�<5>�<`   `   f��<)�<T��<���<_�<�s�<GF�<b��<t��<��<,n�<m��<R��<m��<,n�<��<t��<b��<GF�<�s�<_�<���<T��<)�<`   `   ���<���<}7�<,��<���<�L�<i��<���<���<��<6��<�<H �<�<6��<��<���<���<i��<�L�<���<,��<}7�<���<`   `    ��<��<���<��<���<�X�<e	�<���<�[�<~�<F��<��<���<��<F��<~�<�[�<���<e	�<�X�<���<��<���<��<`   `   �V�<�C�<|�<���<v%�<B�<���<���<�:�<u��<W�<=��<&��<=��<W�<u��<�:�<���<���<B�<v%�<���<|�<�C�<`   `   ԅ�<ce�<��<�l�<��< �<���<!f�<G�<�@�<"l�<C��<��<C��<"l�<�@�<G�<!f�<���< �<��<�l�<��<ce�<`   `   YD�<U�<I��<O��<��<8��<cJ�<��<�P�<���<[��<Q�<���<Q�<[��<���<�P�<��<cJ�<8��<��<N��<I��<U�<`   `   U��<�j�<���<C�<���<�}�<���<��<M4�<7��<�#�<5:�<���<5:�<�#�<7��<M4�<��<���<�}�<���<C�<���<�j�<`   `   ?�<�Q�<���<X��<ז�<���<&�<P��<���<��<rK�<F�<���<F�<rK�<��<���<P��<&�<���<ז�<X��<���<�Q�<`   `   ���<���<M4�<�9�<m��<�<���<Ѝ�<�0�<��<A�<�!�<���<�!�<A�<��<�0�<Ѝ�<���<�<m��<�9�<M4�<���<`   `   ���<l��<m0�<=!�<��<��<�Q�<��<{6�<���<���<���<#X�<���<���<���<{6�<��<�Q�<��<��<=!�<l0�<l��<`   `   -��<�c�<w��<r��<P��<#��<�Z�<��<P��<�q�<Ml�<��<��<��<Ml�<�q�<P��<��<�Z�<#��<O��<r��<v��<�c�<`   `   ���<��<[��<��<���<���<�<D6�<yS�<���<Nz�<��<��<��<Nz�<���<yS�<D6�<�<���<���<��<[��<��<`   `   I��<:a�<���< G�<�u�<#�<�i�<�i�<�U�<�s�<��<1��<���<1��<��<�s�<�U�<�i�<�i�<#�<�u�< G�<���<:a�<`   `   �.�<���<��<<��<���<:K�<Wp�<9A�<��<N��<�2�<kw�<;��<kw�<�2�<N��<��<9A�<Vp�<:K�<���<<��<��<���<`   `   �_�<?�<G!�<��<K��<O$�<�#�<n��<�.�<��<p��<m�<_Y�<m�<p��<��<�.�<n��<�#�<O$�<K��<��<F!�<?�<`   `   `=�<���<[��<�b�<]N�<.��<4��<��<�&�<�{�<sg�<�V�<��<�V�<sg�<�{�<�&�<��<4��<-��<]N�<�b�<[��<���<`   `   ��<@s�<�l�<���<��<K�<��<	�<��<"(�<���<=��<N��<=��<���<"(�<��<	�<��<J�<��<���<�l�<@s�<`   `   ��<��<���<��<���<�>�<?��<n!�<X�<��<���<�m�<֠�<�m�<���<��<X�<m!�<?��<�>�<���<��<���<��<`   `   92�<B��<_��<�0�<u�<Qu�<�7�<zs�<�e�<�r�<7�<C��<�<C��<6�<�r�<�e�<zs�<�7�<Qu�<u�<�0�<^��<B��<`   `   8-�<���<p��<J�<�N�<���<l��<�-�<�T�<���<�`�<�9�<w�<�9�<�`�<���<�T�<�-�<l��<���<�N�<J�<p��<���<`   `   S$�<��<���<ex�<���<�k�<���<�r�<���<{��<H��<���<��<���<H��<{��<���<�r�<���<�k�<���<dx�<���< ��<`   `   �1�<���<<�<��<vN�<Se�<,�<.W�<�a�<cz�<,��<�Q�<f��<�Q�<,��<cz�<�a�<-W�<,�<Se�<vN�<��<<�<���<`   `   `s�<�5�<U��<i��<{K�<���<��<���<���<�9�<A@�<'��<�n�<'��<@@�<�9�<���<���<��<���<{K�<h��<U��<�5�<`   `   ���<h��<-J�<���<u��<��<�f�<_��<�H�<£�<8�<6>�<1��<6>�<8�<£�<�H�<^��<�f�<��<t��<���<-J�<g��<`   `   S��<n��<-n�< �<u��<c��<HF�<�s�<`�<���<U��<*�<g��<*�<T��<���<_�<�s�<GF�<c��<u��<��<-n�<n��<`   `   H �<�<7��<��<���<���<j��<�L�<���<-��<~7�<���<���<���<~7�<-��<���<�L�<j��<���<���<��<7��<�<`   `   ���<��<G��<�<�[�<���<f	�<�X�<���<��<���<��<��<��<���<��<���<�X�<f	�<���<�[�<~�<G��<��<`   `   ��<I��<�V�<_��<���<��<fb�<���<P��<�}�<���<+��<�*�<*��<���<�}�<P��<���<fb�<��<���<_��<�V�<I��<`   `   ���<���<���<�3�<�i�<�s�<�8�<|��<���<N��<��<���<L�<���<��<N��<���<|��<�8�<�s�<�i�<�3�<���<���<`   `   J�<�\�<��<� �<lM�<j�<�N�<���<"�<%�<���<���<��<���<���<%�<"�<���<�N�<j�<lM�<� �<��<�\�<`   `   _��<�S�<j��<O�<!c�<m�<�k�<���<B%�<���<E�<qo�<c�<qo�<E�<���<B%�<���<�k�<m�<!c�<O�<j��<�S�<`   `   ���<Ng�<��<=��<�x�<���<�i�<���<p��<�A�<#�<��<���<��<
#�<�A�<p��<���<�i�<���<�x�<=��<��<Ng�<`   `   ټ�<Us�<9��<���<k�<�a�<�/�<���<�C�<�K�<=��<4c�<C��<4c�<<��<�K�<�C�<���<�/�<�a�<k�<���<9��<Us�<`   `   �k�<�J�<��<���<�"�<7�<��<��<�g�<��<���<2��<�;�<2��<���<��<�g�<��<��<7�<�"�<���<��<�J�<`   `   ���<|��<���<
�<���<�j�<��<�!�<\�<b��<���<(F�<���<(F�<���<b��<\�<�!�<��<�j�<���<
�<���<|��<`   `   �C�<�{�<��<�J�<���<T��<hK�<'E�<E�<�-�<��<N��<(3�<N��<��<�-�<E�<'E�<hK�<T��<���<�J�<��<�{�<`   `   bJ�<λ�<�ޱ<� �<[��<��<���<��<vO�<���<�'�<*�<���<*�<�'�<���<vO�<��<���<��<[��<� �<�ޱ<λ�<`   `   !��<��<��<�Я<���< �<��<��<���<���<���<o�<{��<o�<���<���<���<��<��< �<���<�Я<��<��<`   `   B��<���<�L�<i��<H�<��<��<K��<@��<�p�<���<%W�<�9�<%W�<���<�p�<@��<K��<��<��<H�<i��<�L�<���<`   `   7i�<Р�<��<�v�<��<h�<�o�<��<�
�<F��<:X�<h:�<�3�<h:�<:X�<F��<�
�<��<�o�<h�<��<�v�<��<Р�<`   `   r�<F]�<]S�<�ǔ<KS�<���<�<k-�<$_�<_��<���<���<���<���<���<_��<$_�<k-�<�<���<KS�<�ǔ<]S�<F]�<`   `   Ŭp<��u<�^�<���<�ݚ<�ߨ<�9�<��<E��<�X�<��<p�<0(�<p�<��<�X�<E��<��<�9�<�ߨ<�ݚ<���<�^�<��u<`   `   �Re<�j<��y< w�<3�<���<�R�<�n�<�x�<�H�<2��<D>�<�]�<D>�<2��<�H�<�x�<�n�<�R�<���<3�< w�<��y<�j<`   `   QHa<��f<�u<�@�<qݓ<�#�<��<�»<��<[��<{�<s�<ǒ�<s�<{�<[��<��<�»<��<�#�<qݓ<�@�<�u<��f<`   `   ECe<%Vj<B�x<�1�<2'�<��<9��<�4�<f��<]8�<��<��<���<��<��<]8�<f��<�4�<9��<��<2'�<�1�<B�x<%Vj<`   `   cq<��u<sb�<�?�<��<�~�<�\�<[�<ħ�<���<���<���<2��<���<���<���<ħ�<[�<�\�<�~�<��<�?�<sb�<��u<`   `   c��<H��<.m�<��<�U�</�<܏�<�ƺ<|�<>��< �<<��<��<<��< �<>��<|�<�ƺ<܏�</�<�U�<��<.m�<H��<`   `   �Q�<���<���<�ښ<Mm�<s�<��<�ļ<�2�<K�<?�<�g�<�2�<�g�<?�<K�<�2�<�ļ<��<s�<Mm�<�ښ<���<���<`   `   Q�<W��<�[�<���<6��<dϲ<1��<z��<ð�< ��<߾�<���<I�<���<߾�< ��<ð�<z��<1��<dϲ<6��<���<�[�<W��<`   `   ª�<|��<
g�<+��<���<w��<X��<�#�<���<���<b��<�\�<���<�\�<b��<���<���<�#�<X��<w��<���<+��<
g�<|��<`   `   �~�<�*�<A�<��<�J�<���<��<���<!T�<�1�<���<�x�<\��<�x�<���<�1�<!T�<���<��<���<�J�<��<A�<�*�<`   `   �*�<)��<���<�}�<O��<���<eb�<��<���<^��<�V�<I��<��<I��<�V�<^��<���<��<eb�<���<O��<�}�<���<)��<`   `   L�<���<��<M��<���<{��<�8�<�s�<�i�<�3�<���<���<���<���<���<�3�<�i�<�s�<�8�<{��<���<M��<��<���<`   `   ��<���<���<$�<"�<���<�N�<j�<kM�<� �<��<�\�<I�<�\�<��<� �<kM�<j�<�N�<���<"�<$�<���<���<`   `   b�<po�<E�<���<A%�<���<�k�<l�< c�<O�<i��<�S�<_��<�S�<i��<O�< c�<l�<�k�<���<A%�<���<E�<po�<`   `   ���<��<
#�<�A�<o��<���<�i�<���<�x�<<��<��<Mg�<���<Mg�<��<<��<�x�<���<�i�<���<o��<�A�<
#�<��<`   `   C��<4c�<<��<�K�<�C�<���<�/�<�a�<k�<���<9��<Us�<ؼ�<Ts�<8��<���<k�<�a�<�/�<���<�C�<�K�<<��<4c�<`   `   �;�<1��<���<��<�g�<��<��<7�<�"�<���< ��<�J�<�k�<�J�< ��<���<�"�<6�<��<��<�g�<��<���<1��<`   `   ���<(F�<���<b��<\�<�!�<��<�j�<���<	�<���<{��<���<{��<���<	�<���<�j�<��<�!�<\�<b��<���<(F�<`   `   (3�<M��<��<�-�<E�<'E�<hK�<T��<���<�J�<��<�{�<�C�<�{�<��<�J�<���<T��<gK�<'E�<E�<�-�<��<M��<`   `   ���<*�<�'�<���<vO�<��<���<��<[��<� �<�ޱ<λ�<aJ�<ͻ�<�ޱ<� �<Z��<��<���<��<uO�<���<�'�<*�<`   `   {��<n�<���<���<���<��<��<�<���<�Я<��<��< ��<��<��<�Я<���<�<��<��<���<���<���<n�<`   `   �9�<$W�<���<�p�<@��<K��<��<��<H�<i��<�L�<���<B��<���<�L�<h��<H�<��<��<K��<?��<�p�<���<$W�<`   `   �3�<h:�<:X�<F��<�
�<��<�o�<i�<��<�v�<��<Р�<7i�<Р�<��<�v�<��<h�<o�<��<�
�<F��<:X�<h:�<`   `   ���<���<���<_��<$_�<k-�<�<���<KS�<�ǔ<]S�<F]�<r�<F]�<]S�<�ǔ<KS�<���<�<k-�<#_�<_��<���<���<`   `   0(�<p�<��<�X�<F��<��<�9�<�ߨ<�ݚ<���<�^�<��u<Ƭp<��u<�^�<���<�ݚ<�ߨ<�9�<��<E��<�X�<��<p�<`   `   �]�<D>�<2��<�H�<�x�<�n�<�R�<���<3�< w�<��y<�j<�Re<�j<��y< w�<3�<���<�R�<�n�<�x�<�H�<2��<D>�<`   `   ǒ�< s�<{�<\��<��<�»<��<�#�<rݓ<�@�<�u<��f<RHa<��f<�u<�@�<rݓ<�#�<��<�»<��<\��<{�<s�<`   `   ���<��<��<]8�<g��<�4�<:��<��<2'�<�1�<D�x<&Vj<FCe<&Vj<C�x<�1�<2'�<��<:��<�4�<f��<]8�<��<��<`   `   3��<���<���<���<ŧ�<[�<�\�<�~�<��<�?�<tb�<��u<dq<��u<tb�<�?�<��<�~�<�\�<[�<ħ�<���<���<���<`   `    ��<=��< �<?��<|�<�ƺ<ݏ�</�<�U�<��</m�<I��<c��<I��</m�<��<�U�</�<ݏ�<�ƺ<|�<>��< �<=��<`   `   �2�<�g�<@�<K�<�2�<�ļ<��<s�<Nm�<�ښ<���<���<�Q�<���<���<�ښ<Nm�<s�<��<�ļ<�2�<K�<@�<�g�<`   `   I�<���<��<!��<İ�<{��<2��<fϲ<7��<���<�[�<X��<Q�<X��<�[�<���<7��<eϲ<2��<z��<İ�<!��<߾�<���<`   `   ���<�\�<c��<���<���<�#�<Y��<y��<���<,��<g�<}��<ê�<}��<g�<,��<���<x��<Y��<�#�<���<���<c��<�\�<`   `   ]��<�x�<���<�1�<"T�<���<��<���<�J�<��<B�<�*�<�~�<�*�<B�<��<�J�<���<��<���<"T�<�1�<���<�x�<`   `   #��<�i�<���<A��< ,�<j'�<��<Ȟ�<Wܢ<]h�<5�<�<,��<�<5�<]h�<Vܢ<Ǟ�<��<j'�< ,�<A��<���<�i�<`   `   �x�<�B�<~��<���<���<C��<Va�<�G�<1��<o��<��<�K�<oW�<�K�<��<o��<0��<�G�<Ua�<B��<���<���<~��<�B�<`   `   l��<<��</�<���<�=�<�L�<���<�\�<d�<��<��<Xf�<Qܺ<Xf�<��<��<d�<�\�<���<�L�<�=�<���</�<<��<`   `   ��<�j�<��<��<
��<���<���<���<���<w��<�
�<�x�<8�<�x�<�
�<v��<���<���<��<���<
��<��<��<�j�<`   `   Uӹ<Ѹ�<�E�</�<#_�<��<���<���<�K�<Ҿ�<�|�<���<���<���<�|�<Ҿ�<�K�<���<���<��<#_�<.�<�E�<Ѹ�<`   `   �ް<�+�<�ʵ<�(�<m��<Y�<�>�<���<I��<���< ��<w��<\�<w��< ��<���<I��<���<�>�<Y�<m��<�(�<�ʵ<�+�<`   `   M��<7�<���<��<v��<���<���<�`�<�f�<���</�<���<���<���</�<���<�f�<�`�<���<���<v��<��<���<7�<`   `   n�<���<��<Ѝ�<�v�<��<��<���<���<���<M�<���<�}�<���<M�<���<ߞ�<���<��<��<�v�<Ѝ�<��<���<`   `   �N�<x�<	S�<=��<4!�<ǅ�<8T�<���<3��<rm�<���<�P�<Yn�<�P�<���<rm�<2��<���<8T�<ǅ�<4!�<=��<	S�<w�<`   `   �P<��V<�-i<BR�<�<큤<�h�<�g�<^��<Yg�<i;�<iS�<��<iS�<i;�<Yg�<^��<�g�<�h�<큤<�<BR�<�-i<��V<`   `   20<J�!<��7<��X<bm�<��<��<x��<s��<A�<�1�<P�<��<P�<�1�<A�<s��<x��<��<��<bm�<��X<��7<J�!<`   `   `��;��;��<�*<�Y<�J�<���<:��<4X�<K��<$>�<��<��<��<$>�<K��<4X�<:��<���<�J�<�Y<�*<��<��;`   `   �;o,?;2��;���;t�0<�i<��<v�<c��<H�<���<�<B%�<�<���<H�<c��<v�<��<�i<t�0<���;2��;o,?;`   `   F���(�����:��;d�<6�J<���<)�<w#�<��<C��<��<�,�<��<C��<��<w#�<)�<���<6�J<d�<��;���:�(��`   `   @�q�H{>���2���-;�J�;��0<n�q<}��<H,�<�i�<�"�<���<���<���<�"�<�i�<H,�<}��<n�q<��0<�J�;��-;��2�H{>�`   `   y�������4�-�:�L�;�<<b�a<V��<Y�< Z�<r��<�T�<���<�T�<r��< Z�<Y�<V��<b�a<�<<�L�;-�:�4����`   `   �ƻ�竻�?�	$:�9�;��<��X<�X�<U"�<zG�<a��<�m�<U��<�m�<a��<zG�<U"�<�X�<��X<��<�9�;	$:�?��竻`   `   !��������V��_w:${�;�<��W<�Ј<{۠<x�<'|�<��<L��<��<'|�<x�<{۠<�Ј<��W<�<${�;�_w:�V�����`   `   'to���?���_��w;�p�;T�!<q^<O7�<��<��<�T�<r��<i��<r��<�T�<��<��<O7�<q^<T�!<�p�;�w;��_���?�`   `   �wc���j����:r��;��;�6<�ml<![�<��<�3�<�C�<���<���<���<�C�<�3�<��<![�<�ml<�6<��;r��;���:��j�`   `   ��+;��O;,��;J��;!^!<��Q<l�<�ʔ<��<⫳<�H�<���<|��<���<�H�<⫳<��<�ʔ<l�<��Q<!^!<J��;,��;��O;`   `   )��;�; <�%<�xJ<��q<���<I�<�#�<O�<�D�<>	�<_��<>	�<�D�<O�<�#�<I�<���<��q<�xJ<�%< <�;`   `   ��*<�P0<�E@<�SX<�]u<��<�ט<�<
�<
��<s �<N��<W�<N��<s �<	��<
�<�<�ט<��<�]u<�SX<�E@<�P0<`   `   h<))l<��w<aބ<���<��<	ʥ<�a�<�S�<��<��<���<��<���<��<��<�S�<�a�<	ʥ<��<���<aބ<��w<))l<`   `   +��<�<5�<\h�<Uܢ<ƞ�<��<i'�<�+�<@��<���<�i�<#��<�i�<���<@��<�+�<i'�<��<ƞ�<Uܢ<\h�<5�<�<`   `   nW�<�K�< ��<n��</��<�G�<Ta�<B��<���<���<}��<�B�<�x�<�B�<}��<���<���<B��<Ta�<�G�</��<n��< ��<�K�<`   `   Pܺ<Wf�<��<��<d�<�\�<���<�L�<�=�<���</�<;��<k��<;��</�<���<�=�<�L�<���<�\�<d�<��<��<Wf�<`   `   8�<�x�<�
�<v��<���<���<��<���<	��<��<��<�j�<��<�j�<��<��<	��<���<��<���<���<u��<�
�<�x�<`   `   ���<���<�|�<Ѿ�<�K�<���<���<~��<"_�<.�<�E�<и�<Tӹ<и�<�E�<.�<"_�<~��<���<���<�K�<Ѿ�<�|�<���<`   `   [�<v��<��<���<H��<���<�>�<X�<l��<�(�<�ʵ<�+�<�ް<�+�<�ʵ<�(�<l��<X�<�>�<���<H��<���<��<v��<`   `   ��<���<.�<���<�f�<�`�<���<���<u��<��<���<7�<M��<7�<���<��<u��<���<���<�`�<�f�<���<.�<���<`   `   �}�<���<L�<���<ߞ�<���<��<��<�v�<ύ�<��<���<n�<���<��<ύ�<�v�<��<��<���<ߞ�<���<L�<���<`   `   Xn�<�P�<���<rm�<2��<���<7T�<ǅ�<4!�<=��<S�<w�<�N�<w�<S�<<��<4!�<ǅ�<7T�<���<2��<qm�<���<�P�<`   `   ��<iS�<i;�<Yg�<^��<�g�<�h�<큤<�<AR�<�-i<��V<�P<��V<�-i<AR�<�<쁤<�h�<�g�<^��<Xg�<i;�<iS�<`   `   ��<P�<�1�<A�<s��<x��<��<��<am�<��X<��7<I�!<10<I�!<��7<��X<am�<��<��<x��<s��<A�<�1�<P�<`   `   ��<��<$>�<J��<4X�<:��<���<�J�<�Y<�*<��<
��;^��;	��;��<�*<�Y<�J�<���<:��<4X�<J��<$>�<��<`   `   B%�<�<���<H�<d��<v�<��<�i<t�0<���;2��;n,?;�;m,?;1��;���;s�0<�i<��<v�<c��<G�<���<�<`   `   �,�<��<C��<��<x#�<)�<���<6�J<e�<��;���:�(��H���(�����:��;d�<5�J<���<)�<w#�<��<C��<��<`   `   ���<���<�"�<�i�<H,�<}��<o�q<��0<�J�;��-;��2�G{>�@�q�H{>���2���-;�J�;��0<n�q<|��<H,�<�i�<�"�<���<`   `   ���<�T�<s��< Z�<Y�<V��<c�a<�<<�L�;-�:�4����x�������4�-�:�L�;�<<b�a<V��<Y�< Z�<s��<�T�<`   `   V��<�m�<a��<{G�<V"�<�X�<��X<��<�9�;$:�?��竻�ƻ�竻�?�$:�9�;��<��X<�X�<U"�<zG�<a��<�m�<`   `   L��<��<(|�<x�<|۠<�Ј<��W<�<'{�;`w:�V�������������V�`w:%{�;�<��W<�Ј<{۠<x�<(|�<��<`   `   j��<s��<�T�<��<��<P7�<q^<V�!<�p�;�w;��_��?�"to��?���_��w;�p�;U�!<q^<P7�<��<��<�T�<s��<`   `   ���<���<�C�<�3�<��<"[�<�ml<�6<��;v��;���:2�j��wc�D�j����:t��;��;�6<�ml<![�<��<�3�<�C�<���<`   `   }��<���<�H�<䫳<��<�ʔ<m�<��Q<#^!<O��;0��;��O;�+;��O;/��;M��;"^!<��Q<m�<�ʔ<��<㫳<�H�<���<`   `   `��<?	�<�D�<�O�<�#�<K�<���<��q<�xJ<�%<<�;.��;�;<�%<�xJ<��q<���<J�<�#�<O�<�D�<?	�<`   `   X�<O��<t �<��<�<�<�ט<��<�]u<�SX<�E@<�P0< �*<�P0<�E@<�SX<�]u<��<�ט<�<�<
��<s �<O��<`   `   ��<���<��<��<�S�<�a�<
ʥ<��<���<bބ<��w<+)l<h<+)l<��w<bބ<���<��<
ʥ<�a�<�S�<��<��<���<`   `   Ժ<ŋ�<���<��<D��<LX�<�;�<�q<�+M<�*<b�<y��;���;y��;b�<�*<�+M<�q<�;�<LX�<C��<��<���<ŋ�<`   `   ���<��<�<&��<O��<g��<ǂ�<��<S�<�x<~e<�W<�)S<�W<~e<�x<R�<��<ǂ�<g��<O��<%��<�<��<`   `   ٷ�<�<ꌵ<��<_
�<+ر<r(�<���<���<�-�<�[�<�M�<�Ӑ<�M�<�[�<�-�<���<���<q(�<+ر<_
�<��<ꌵ<ﰵ<`   `   0í<�a�<�#�<���<�j�<ޙ�<;��</e�<:۶<�<�<��<1f�<��<�<�<:۶<.e�<:��<ޙ�<�j�<���<�#�<�a�<`   `   ���<��<ȥ<Oh�<t�<nY�< ۽<Y��<���< ��<I%�<��<�	�<��<I%�< ��<���<Y��< ۽<nY�<t�<Oh�<ȥ<��<`   `   ^4�<�P�<V�<�F�<B֨<���<0��<K��<�X�<r��<]��<�H�<O��<�H�<]��<q��<�X�<K��<0��<���<B֨<�F�<V�<�P�<`   `   	�d<��j<t�{<u�<��<)�<��<7��<���<Tx�<���<���<I��<���<���<Tx�<���<7��<��<)�<��<u�<t�{<��j<`   `   Ѷ<R�&<�=<��^<���<<��<��<AX�<ī�<���<t.�<Y��<[*�<Y��<s.�<���<ī�<AX�<��<<��<���<��^<�=<R�&<`   `   �;vܢ;�v�;��<=�M<�N�<�p�<�r�<�T�<)��<���<F��<���<F��<���<)��<�T�<�r�<�p�<�N�<=�M<��<�v�;vܢ;`   `   �\������a:O�;�8<�AM<��<}��<�s�<���<���<
�<���<
�<���<���<�s�<}��<��<�AM<�8<O�;�a:����`   `   6��D�ķ��v���[<c;E}<�*^<ӟ�< �<LN�<���<���<���<���<���<KN�< �<ӟ�<�*^<E}<Z<c;w���ķ���D�`   `   �7��P�����N�xT��������;)<��}<���<�+�<L��<Q�<��<Q�<L��<�+�<���<��}<)<���;���xT����N�P���`   `   � ͼS���*���0d��!���b9�i�;=U<��<L�<�x�<Y��<���<Y��<�x�<L�<��<=U<�i�;��b9�!�0d�*���S���`   `   �z�V��b�׼�t��HB���s�Q��;��.<�G�<:~�<��<��<:�<��<��<:~�<�G�<��.<Q��;��s�HB��t��b�׼V��`   `   ��j������jȼ����>廅q�:��<�o<��<7�<v��<��<v��<7�<��<�o<��<�q�:�>廘���jȼ���j��`   `   �!-�u�%����?�⼖���� �=U��W�;��Z<gA�<��<V��<~��<V��<��<gA�<��Z<�W�;>U�� �����?�⼒��u�%�`   `   ��2��D+����'���ۡ��8)�M������;|�M<�7�<�U�<��<X(�<��<�U�<�7�<|�M<���;M����8)��ۡ�'�켟���D+�`   `   L!-���%�$>�aC��֜�[�#�m���c�;tI<0�<Up�<hմ<$ع<hմ<Up�<0�<tI<c�;m���[�#��֜�aC�$>���%�`   `   >��� �����4ͼ� �����O
��y�;7�L<r�<2��<�<�ڶ<�<2��<r�<7�L<y�;P
������ ���4ͼ���� �`   `   ���,-���vټ 4����V�} ��w�:2�<�DX<��<躣<^��<8S�<^��<躣<��<�DX<2�<w�:} ����V� 4���vټ,-��`   `   I�ȼ�������n���#9�r��;�P <�j<Zޑ<�ѥ<�p�<{<�<�p�<�ѥ<Zޑ<�j<�P <r��;$9����n�������`   `   �p���x�,"J����`
E�!�;��;D�C<Oˀ<���<�l�<�4�<]i�<�4�<�l�<���<Oˀ<D�C<��;!�;`
E����,"J��x�`   `   G ���D)���Oź��";@�;��/<vRj<`��<���<�<��<GG�<��<�<���<`��<vRj<��/<@�;��";�OźD)����`   `   ]��7��:�3;�ț;>,�;��2<Pod<�#�<�N�<�d�<�K�<��<�
�<��<�K�<�d�<�N�<�#�<Pod<��2<>,�;�ț;�3;��:`   `   ���;t��;_�<�*<�+M<�q<�;�<KX�<B��<��<��<ċ�<Ժ<ċ�<��<��<B��<KX�<�;�<�q<�+M<�*<_�<t��;`   `   �)S<�W<{e<�x<Q�<��<Ƃ�<f��<N��<$��<�<��<���<��<�<$��<N��<f��<Ƃ�<��<Q�<�x<{e<�W<`   `   �Ӑ<�M�<�[�<�-�<���<���<p(�<*ر<^
�<��<錵<ﰵ<ط�<ﰵ<錵<��<^
�<*ر<p(�<���<���<�-�<�[�<�M�<`   `   0f�<��<�<�<9۶<-e�<:��<ݙ�<�j�<���<�#�<�a�</í<�a�<�#�<���<�j�<ݙ�<9��<-e�<9۶<�<�<��<`   `   �	�<��<H%�<��<���<X��<۽<mY�<s�<Nh�<ȥ<��<���<��<ȥ<Nh�<s�<mY�<۽<X��<���<��<G%�<��<`   `   N��<�H�<\��<q��<�X�<J��</��<���<B֨<�F�<V�<�P�<]4�<�P�<V�<�F�<A֨<���</��<J��<�X�<p��<\��<�H�<`   `   H��<���<���<Sx�<���<6��<��<)�<��<u�<s�{<��j<�d<��j<s�{<u�<��<)�<��<6��<���<Sx�<���<���<`   `   Z*�<X��<s.�<���<ë�<@X�<��<;��<���<��^<�=<P�&<϶<P�&<�=<��^<���<;��<��<@X�<ë�<���<s.�<X��<`   `   ���<F��<���<(��<�T�<�r�<�p�<�N�<<�M<��<�v�;tܢ;;sܢ;�v�;��<<�M<�N�<�p�<�r�<�T�<(��<���<F��<`   `   ���<
�<���<���<�s�<|��<��<�AM<�8<M�;�a:�����\������a:L�;�8<�AM<��<|��<�s�<��<���<
�<`   `   ���<���<���<KN�<�߯<ӟ�<�*^<E}<X<c;}���Ʒ���D�7��D�Ƿ������U<c;D}<�*^<ҟ�<�߯<KN�<���<���<`   `   ��<Q�<L��<�+�<���<��}<)<���;���yT����N�Q����7��Q�����N�zT��������;)<��}<���<�+�<L��<Q�<`   `   ���<Y��<�x�<L�<��<=U<�i�;��b9�!�0d�*���S���� ͼT���+���1d��!廮�b9�i�;<U<��<L�<�x�<X��<`   `   :�<��<��<:~�<�G�<��.<R��;��s�HB��t��b�׼V���z�V��c�׼�t��HB���s�O��;��.<�G�<:~�<��<��<`   `   ��<v��<7�<���<�o<��<�q�:�>廘���jȼ��j����j������jȼ����>廁q�:��<�o<��<7�<v��<`   `   ~��<W��<��<hA�<��Z<�W�;+U�� �����>�⼒��u�%��!-�u�%����?�⼖���� �?U��W�;��Z<hA�<��<W��<`   `   Y(�<��<�U�<�7�<~�M<���;A����8)��ۡ�'�켞���D+���2��D+����'���ۡ��8)�K������;|�M<�7�<�U�<��<`   `   %ع<iմ<Vp�<1�<vI<c�;^���Y�#��֜�`C�#>���%�L!-���%�#>�aC��֜�Z�#�i���c�;uI<0�<Vp�<iմ<`   `   �ڶ<�<3��<s�<9�L<}�;
������ ���4ͼ���� �=��� �����4ͼ� �����6
��{�;8�L<s�<3��<�<`   `   9S�<_��<꺣<��<�DX<4�<(w�:x ����V��3���vټ+-�����+-���vټ 4����V�z ��w�:3�<�DX<��<麣<_��<`   `   |<�<�p�<�ѥ<[ޑ<�j<�P <w��;9����n�������H�ȼ�������n���9�u��;�P <�j<Zޑ<�ѥ<�p�<`   `   ^i�<�4�<�l�<���<Pˀ<G�C<#��;,�;U
E����)"J��x��p���x�*"J����Z
E�(�;!��;E�C<Pˀ<���<�l�<�4�<`   `   HG�<��<�<���<a��<yRj<��/<@�;��";�Oź?)����E ���@)���Oź��";@�;��/<wRj<a��<���<�<��<`   `   �
�<��<�K�<�d�<�N�<�#�<Sod<��2<D,�;ɛ;�3;��:���7��:�3; ɛ;C,�;��2<Rod<�#�<�N�<�d�<�K�<��<`   `   ���<獨<�<�;�<���<�Q<��<:�;tx�9�=z�*���� ���.��� �+���=z�Wx�9:�;��<�Q<���<�;�<�<獨<`   `   �<׊�<g^�<���<��<w��<!^<
�1<�z<1b�;�&,;�\�:^�9�\�:�&,;0b�;�z<	�1< ^<v��<��<���<g^�<׊�<`   `   k�<�#�<�!�<���<��<���<5��<�Z}<b<	HF<I(.<r�<�<r�<I(.<	HF<b<�Z}<5��<���<��<���<�!�<�#�<`   `   ���<_V�<Ď�<���<�z�<K �<*��<��<���<Q��<g�<Cʄ<�P�<Cʄ<g�<Q��<���<��<*��<K �<�z�<���<Ď�<_V�<`   `   G�s<k�w<���<��<�ٓ<�;�<Y�<��<�<�?�<���<�<T��<�<���<�?�<<��<Y�<�;�<�ٓ<��<���<k�w<`   `   ��*<�I1<̧D<3�a<��<&X�<J1�<�4�<D�<_t�<��<��<yj�<��<��<_t�<D�<�4�<J1�<&X�<��<3�a<̧D<�I1<`   `   !#�;jD�;���;G<��H<�}<W��<g��<,��<f��<�[�<=(�<���<=(�<�[�<e��<,��<g��<W��<�}<��H<G<���;jD�;`   `   �.�O���E�G;;'��;�><4.�<#d�<��<�_�<��<rd�<���<rd�<��<�_�<��<"d�<3.�<�><'��;G;;��E�/�O�`   `   ��k�\!Y��n$�@X����:h�;��F<<�<��<Q�<.E�<�@�<؀�<�@�<.E�<P�<��<<�<��F<h�;��:@X���n$�\!Y�`   `   �|ܼjwм�[��̷v�8���=�8���;۪`<�ܚ<�#�<�Y�<�-�<9X�<�-�<�Y�<�#�<�ܚ<ڪ`<���;$�88���̷v��[��jwм`   `   Վ)���!�fL�B ؼ}���W���:vO<��<��<��<�a�<ч�<�a�<��<��<��<uO<���:W�}���B ؼfL���!�`   `   ҄j�~a��GF�i���B߼�}����	�;�BT<=�<��<+��<*�<+��<��<<�<�BT<�	�;���}��B߼i���GF�~a�`   `   V���Ґ�J���)�Q���f�����-��!:�p<G��<L!�<�!�<K�<�!�<L!�<G��<�p<�!:��-�f�����)�Q�J���Ґ�`   `   ֱ������p��������A�� �Ҝ��Gr��D�;��h<>'�<�ݷ<~�<�ݷ<>'�<��h<�D�;Hr�Ҝ��� ���A������p�����`   `   �sϽȽ�Q��E͔��mb�X������)�\z;=6G<�8�<��<Hյ<��<�8�<=6G<\z;�)񻁛��X��mb�E͔��Q��Ƚ`   `   ���E�ؽ½����x��,���ʼjd$��]�:fs,<@D�<%��<}Ŭ<%��<@D�<fs,<�]�:jd$���ʼ�,���x���½E�ؽ`   `   ����޽|Ƚ���GÀ��3�
/ؼ3z;�c:<�<�?~<!�<�F�< �<�?~<;�<c:3z;�
/ؼ�3�GÀ����|Ƚ��޽`   `   ��ཎ�ؽý�����{�C0�Sռ�y;�N�z9�<9�t<&��<)ܟ<&��<9�t<�<L�z9�y;�SռC0���{����ý��ؽ`   `   �=Ͻ�Ƚ���E����9h�"�l¼�$�qbt:�;<8�r<��<�֜<��<8�r<�;<qbt:�$�l¼"��9h�E�������Ƚ`   `   �������(������!I�-�
�/1��+�8$;��#<��w<�\�<�V�<�\�<��w<��#<8$;+�/1��-�
��!I����(������`   `   �ޔ�ꠏ�р�*�U��"�m�ټ�!l���z�J�;R�9<i��<�'�<5(�<�'�<i��<R�9<J�;��z��!l�m�ټ�"�*�U�р�ꠏ�`   `   ��d��K\��rD��� �X��於��	�_�9�Z�;�jU<�ŉ<қ<��<қ<�ŉ<�jU<�Z�;^�9��	��於X���� ��rD��K\�`   `   `� ��A�8��wؼY喼�%��_��m�;��+<t�s<ݺ�<�/�<��<�/�<ݺ�<t�s<��+<�m�;�_��%�Y喼wؼ8���A�`   `   Elļ����J?��� l�h�	�}��_�x;��<�yZ<�J�<V	�<P�<Iv�<P�<V	�<�J�<�yZ<��<_�x;}��h�	�� l�J?������`   `   ��.��� �0���=z�x�9:�;��<�Q<���<�;�<
�<捨<���<捨<
�<�;�<���<�Q<��<:�;x�9�=z�0���� �`   `    �9p\�:w&,;+b�;�z<�1<^<u��<��<���<f^�<֊�<�<֊�<f^�<���<��<u��<^<�1<�z<+b�;w&,;p\�:`   `   	�<o�<F(.<HF<�b<�Z}<4��<���<��<���<�!�<�#�<k�<�#�<�!�<���<��<���<4��<�Z}<�b<HF<F(.<o�<`   `   �P�<Bʄ<f�<P��<���<��<)��<J �<�z�<���<Î�<^V�<���<^V�<Î�<���<�z�<J �<)��<��<���<P��<f�<Bʄ<`   `   S��<�<���<�?�<<��<X�<�;�<�ٓ<��<���<i�w<E�s<i�w<���<��<�ٓ<�;�<X�<��<<�?�<���<�<`   `   wj�<��<��<^t�<C�<�4�<I1�<%X�<��<2�a<ʧD<�I1<��*<�I1<ʧD<1�a<��<%X�<I1�<�4�<C�<^t�<��<��<`   `   ���<=(�<�[�<e��<+��<f��<V��<�}<��H<E<���;gD�;#�;gD�;���;E<��H<�}<V��<f��<+��<d��<�[�<<(�<`   `   ���<qd�<��<�_�<��<"d�<3.�<�><$��;G;;�E�5�O��6�O��E�G;;#��;�><3.�<"d�<��<�_�<��<qd�<`   `   ׀�<�@�<-E�<P�<��<;�<��F<h�;��:BX���n$�]!Y���k�]!Y��n$�CX����:h�;��F<;�<��<P�<-E�<�@�<`   `   8X�<�-�<�Y�<#�<�ܚ<ڪ`<���;��8:���ͷv��[��kwм�|ܼkwм�[��ͷv�;���^�8���;٪`<�ܚ<#�<�Y�<�-�<`   `   ч�<�a�<��<��<��<uO<���: W�}���B ؼfL���!�֎)���!�gL�B ؼ~���"W���:tO<��<��<��<�a�<`   `   *�<+��<��<<�<�BT<�	�;���}��B߼i���GF�~a�ӄj�~a��GF�i���B߼�}����	�;�BT<<�<��<+��<`   `   K�<�!�<L!�<G��<�p<�!:��-�f�����)�Q�J���Ґ�V���Ґ�J���)�Q���g�����-��!:�p<G��<L!�<�!�<`   `   ~�<�ݷ<>'�< �h<�D�;Er�Ҝ��� ���A������p�����ֱ������p��������A�� �Ӝ��Jr��D�;��h<>'�<�ݷ<`   `   Hյ<��<�8�<>6G<_z;�)񻀛��X��mb�E͔��Q��Ƚ�sϽȽ�Q��E͔��mb�X������)�[z;=6G<�8�<��<`   `   ~Ŭ<%��<@D�<gs,<�]�:id$���ʼ�,���x���½E�ؽ���E�ؽ½����x��,���ʼjd$��]�:fs,<@D�<%��<`   `   �F�<!�<�?~<=�< c:2z;�	/ؼ�3�GÀ����|Ƚ��޽����޽|Ƚ���GÀ��3�	/ؼ3z;�c:<�<�?~<!�<`   `   )ܟ<'��<;�t<�<ɒz9�y;�RռC0���{����ý��ؽ��ཎ�ؽý�����{�C0�Sռ�y;�t�z9�<:�t<'��<`   `   �֜<��<:�r<�;<�bt:�$�k¼"��9h�D�������Ƚ�=Ͻ�Ƚ���D����9h�"�l¼�$�bt:�;<:�r<��<`   `   �V�<�\�<��w<��#<8$;&�-1��,�
��!I����'�������������'������!I�,�
�.1��)�8$;��#<��w<�\�<`   `   6(�<�'�<j��<T�9<P�;��z��!l�l�ټ�"�)�U�р�頏��ޔ�頏�р�)�U��"�l�ټ�!l���z�M�;S�9<j��<�'�<`   `   ��<қ<�ŉ<�jU<�Z�;��9��	��於V���� ��rD��K\���d��K\��rD��� �W��於��	���9�Z�;�jU<�ŉ<қ<`   `   ��<�/�<޺�<w�s<��+<�m�;�_��%�W喼vؼ8���A�_� ��A�8��vؼX喼�%��_��m�;��+<v�s<޺�<�/�<`   `   Jv�<Q�<W	�<�J�<zZ<��<l�x;p��e�	�� l�I?������Dlļ����I?��� l�f�	�u��g�x;��<zZ<�J�<W	�<Q�<`   `   `��<$Ґ<���<�Z</�<9Ђ;��)���&�@�����ռ��\�z���\����ռA�����&���)�7Ђ;.�<
�Z<���<$Ґ<`   `   �f�<��<���<{Tt<��K<C <3y�;>}��4���|.���v�듼����듼��v��|.�4���}��1y�;B <��K<zTt<���<��<`   `   H��<��<ˮ�<%�y<r�h<#O<�+<���;3d�;-Һ:Hw��PL�6�v�QL�Kw��(Һ:1d�;���;�+<#O<q�h<$�y<ˮ�<��<`   `   D%V<7gX<7Z^<~�e<@�k<�{l<d�e<WGW<�B<g�)<�<iS<���;iS<�<g�)<�B<VGW<c�e<�{l<?�k<}�e<6Z^<7gX<`   `   ջ<B�<�4<�2<�SO<yZj<�r<�!�<5r�<���<���<6��<�ڂ<6��<���<���<5r�<�!�<�r<yZj<�SO<��2<�4<B�<`   `   �K9�^:v�1;9�;V�<BPF<@Jw<f�<EƝ<�5�<�ʬ<C��<�n�<B��<�ʬ<�5�<EƝ<f�<?Jw<APF<V�<9�;u�1;�^:`   `   :�.�����߻��'��A#;P��;V�M<i��<��<�k�<�-�<1N�<���<1N�<�-�<�k�<��<i��<V�M<P��;�A#;��'���߻��`   `   ��μ�.ü󾡼(�_��ӻ�)�:��<f�e<�y�<��<m�<���<�/�<���<m�<��<�y�<e�e<��<�)�:�ӻ(�_�󾡼�.ü`   `   V4��2,�w4�R �/j��&�n|�:"�<�؅<馮<�n�<�W�<�{�<�W�<�n�<馮<�؅<"�<l|�:&�/j��R �w4��2,�`   `   �����'��8�i�m<�D~��ូlf�#�;�9N<�R�<N��<�X�<p�<�X�<N��<�R�<�9N<"�;lfỬូD~�m<�8�i��'��`   `   ����v�� o���ሽ��L�V�������H��� <C2�<���<Ñ�<��<Ñ�<���<C2�<�� <��H����V����L��ሽ o���v��`   `   � ��&���ݽ_��D���l�A���781��$;lK<�]�<һ<��<һ<�]�<lK<�$;781���l�A�D���_���ݽ�&��`   `   �� ��B����������T�����꙼<<H�y�<�<�ת<�̶<�ת<�<y�<<<H��꙼����T����������B�`   `    @�7�9���&����Nڽ����3rI�w�׼0	���;D�_<�Z�<�ަ<�Z�<D�_<��;0	�w�׼3rI������Nڽ����&�7�9�`   `   �]Z��R���=�ы�O���̼���cm�l��PT��e�:�)7<���<���<���<�)7<�e�:PT�l���cm�̼��O���ы���=��R�`   `   ��k���c��NM���,��{��RŽ?������Ӆ��#���
<u�u<E��<u�u<�
<�#���Ӆ����?���RŽ�{���,��NM���c�`   `   �/r���i���R��1�+��81̽m∽��!��E����/����;S�`<@7�<S�`<���;��/��E����!�m∽81̽+���1���R���i�`   `   ��k�d�c�̫M��m-�t���jȽ)ꆽ�� �TŖ�iP�WJ�;��S<%�r<��S<WJ�;iP�TŖ��� �)ꆽ�jȽt���m-�̫M�d�c�`   `   �0Z���R�Fw>�@� ���������7{�]8�i��¬&����;�P<�m<�P<���;¬&�i��]8��7{��������@� �Fw>���R�`   `   m�?��39�;t'����.�߽=�� >\��� ��Tc���c��.<�TU<�vp<�TU<�.<��c��Tc��� � >\�=��.�߽���;t'��39�`   `   ���{X�+�� S�g���OF��Tp4� ̼��iO�:)y<�xb<Pz<�xb<)y<iO�:�� ̼Tp4�OF��g��� S�+��{X�`   `   ����'��nRܽ��V+���	S�������U��
	�;,27<3�t<&X�<3�t<,27<
	�;�U��������	S�V+����nRܽ'��`   `   ����մ�T#��D����pT��\�")������9�<��V<��<��<��<��V<�<�9���")���\��pT�D���T#���մ�`   `   �퀽F�x���^��C8�U�
�rٷ���?�<����;��2<�\s<CN�<!\�<CN�<�\s<��2<��;<����?�rٷ�U�
��C8���^�F�x�`   `   {���\����ռB�����&���)�3Ђ;,�<�Z<���<#Ґ<_��<#Ґ<���<�Z<,�<3Ђ;��)���&�B�����ռ��\�`   `   ����듼��v��|.� 4���~��-y�;@ <��K<xTt<���<��<�f�<��<���<xTt<��K<@ <-y�;�~�� 4���|.���v�듼`   `   B�v�]L�`w��Һ:-d�;���;�+<#O<o�h<"�y<ʮ�<��<G��<��<ʮ�<"�y<o�h<#O<�+<���;,d�;Һ:aw��]L�`   `   ڎ�;fS<�<d�)<�B<TGW<a�e<�{l<=�k<{�e<4Z^<5gX<B%V<5gX<4Z^<{�e<=�k<�{l<a�e<TGW<�B<d�)<�<fS<`   `   �ڂ<5��<���<���<4r�<�!�<�r<wZj<�SO<�2<�4<@�<ӻ<@�<�4<�2<�SO<wZj<�r<�!�<4r�<���<���<5��<`   `   �n�<A��<�ʬ<�5�<DƝ<f�<=Jw<?PF<T�<9�;n�1;��^:��K9��^:m�1;9�;T�<?PF<=Jw<f�<DƝ<�5�<�ʬ<A��<`   `   ���<0N�<�-�<�k�<��<h��<T�M<M��;�A#;��'���߻��<�.�����߻��'��A#;L��;T�M<h��<��<�k�<�-�<0N�<`   `   �/�<���<l�<��<�y�<d�e<��<�)�:�ӻ)�_�󾡼�.ü��μ�.ü����*�_�	�ӻ�)�:��<c�e<�y�<��<l�<���<`   `   �{�<�W�<�n�<覮<�؅<!�<c|�:'�0j��S �w4��2,�V4��2,�w4�S �0j��(�^|�: �<�؅<覮<�n�<�W�<`   `   o�<�X�<M��<�R�<�9N<!�;nfỬូE~�m<�9�i��'�������'��9�i�m<�E~��ូof��;�9N<�R�<M��<�X�<`   `   ��<Ñ�<���<C2�<�� <��H����V����L��ሽ o���v�������v��!o���ሽ��L�V�������H��� <C2�<���<Ñ�<`   `   ��<һ<�]�<lK<�$;881���l�A�D���_���ݽ�&��� ��&���ݽ_��D���l�A���981�
�$;kK<�]�<һ<`   `   �̶<�ת<�<y�<<<H��꙼����T����������B��� ��B����������T�����꙼@<H�x�<�<�ת<`   `   �ަ<�Z�<E�_<��;/	�w�׼3rI������Nڽ����&�7�9� @�7�9���&����Nڽ����3rI�x�׼0	���;D�_<�Z�<`   `   ���<���<�)7<�e�:OT�l���cm�̼��O���ы���=��R��]Z��R���=�ы�O���̼���cm�l��PT��e�:�)7<���<`   `   E��<v�u<�
<�#���Ӆ����?���RŽ�{���,��NM���c���k���c��NM���,��{��RŽ?������Ӆ��#���
<v�u<`   `   @7�<T�`<���;��/��E����!�m∽81̽+���1���R���i��/r���i���R��1�+��81̽m∽��!��E����/����;T�`<`   `   '�r<��S<[J�;iP�SŖ��� �)ꆽ�jȽt���m-�˫M�d�c���k�d�c�˫M��m-�t���jȽ)ꆽ�� �TŖ�	iP�YJ�;��S<`   `   �m<�P<���;��&�i��]8��7{��������@� �Fw>���R��0Z���R�Fw>�@� ���������7{�]8�i����&����;�P<`   `   �vp<�TU<�.<��c��Tc��� �>\�=��.�߽���;t'��39�m�?��39�;t'����.�߽=�� >\��� ��Tc���c��.<�TU<`   `   Pz<�xb<,y<O�:�� ̼Tp4�OF��f��� S�+��{X����{X�+�� S�g���OF��Tp4� ̼��uO�:+y<�xb<`   `   'X�<6�t</27<	�;�U��첎�����	S�V+����nRܽ'�����'��nRܽ��V+���	S����첎��U��	�;.27<5�t<`   `   ��< 	�<��V<�<t�9���!)���\��pT�D���T#���մ�����մ�T#��D����pT��\�!)�����J�9�<��V< 	�<`   `   "\�<DN�<�\s<��2<��;/����?�pٷ�T�
��C8���^�E�x��퀽E�x���^��C8�T�
�qٷ���?�5����;��2<�\s<DN�<`   `   �wo<b<�8<���;��9�G
�F�8��FZ<���s�$p��]o�����]o��$p����s�FZ<�8��G򞼈G
���9���;�8<b<`   `   ]�c<'F\<^�C<<7��;�!�����oC���˼�)
��1)�<,>��E�<,>��1)��)
��˼oC�����"��5��;<^�C<&F\<`   `   �!;<�8<Ѭ0<��<
�<^m�;l)�:f�\����>f��ؘ��i���x���i���ؘ��>f�	��j�\�d)�:\m�;	�<��<Ь0<�8<`   `   ,e�;w��;.,�;��;�<O� <O�;2��;�:;@�9	�	�CIu��덻DIu��	��?�9�:;0��;�N�;N� <�<��;-,�;w��;`   `   ~캇���o۶9��,;˩;� �;k< �&<��)<f�#<�<�<�d<�<�<f�#<��)<��&<~k<� �;˩;��,;c۶9����`   `   �j�@�Y���*�V�ɻ�!���|;!�<�A<<�j<���<�̉<*�<��<*�<�̉<���<;�j<�A< �<�|;�!��W�ɻ��*�A�Y�`   `   v������k�ռ	����;��[���;d�)<#�y<�<��<�0�<5b�<�0�<��<�<#�y<c�)<��;�[��;�	���k�ռ����`   `   �8h���^��]C�P���ּk�bS[�D��;��\<^\�<�X�<S=�<E��<S=�<�X�<]\�<��\<C��;cS[�k��ּP���]C���^�`   `   65��TW��M ����~�a3<��\𼆸e��Q{��h<	
�<qS�<�a�<'�<�a�<qS�<	
�<�h<�Q{���e��\�a3<���~�M ��TW��`   `   x���9 ���T���G��O�E��{�s�)�L�_;m
^<~ܦ<l��<��<l��<~ܦ<m
^<K�_;s�)��{�O�E�G��T������9 �`   `   ��7�^\1�;`�A%�>�ͽ~Y���5��������<8�<�}�<j��<�}�<8�<�<�������5�~Y��>�ͽA%�;`�^\1�`   `   �9r�<�i�?R��#0�3	��=Ž9���E���P���H;��^<�z�<�a�<�z�<��^<��H;��P��E�9���=Ž3	��#0�?R�<�i�`   `   .����(���B��(�]�1-�<U��.�� |C��뱼�B��<7D�<V�<7D�<�<�B��뱼 |C�.��<U��1-�(�]��B���(��`   `   �H���°�᭞�C؄���O�cs���˽��v�\\��R�����;��Z<��<��Z<���;R��\\����v���˽cs���O�C؄�᭞��°�`   `    �Ѿ�ʾ�7��������l�b0-�:,�]P���`��e���:��*<F�Y<��*<��:�e��`�]P��:,�b0-���l������7���ʾ`   `   z���U۾ �ľ4C��q��� <��o ��Π�w0�����κ��!	<�M4<!	<κ������w0��Π��o �� <�q��4C�� �ľ�U۾`   `   ����~�1ʾ����C���(B�y#�&��6<��t����W����;��<���;��W��t��6<�&��y#��(B�C������1ʾ�~�`   `   0�㾗e۾K�ľCԤ��O��"c>��as���<�P}��������;"w<���;���P}���<�as���"c>��O��CԤ�K�ľ�e۾`   `   �Ѿ�ʾ����ᅘ�Np�_1��������b0��w���[o��;X�<�;�[o��w��b0��������_1�Np�ᅘ������ʾ`   `   "Զ���,��W����S����>ٽ���̧�bޅ�n	� �;��<	 �;n	�bޅ�̧�����>ٽ���S�W���,����`   `   Í��;u��mF��]�_�`c1�'���=����e�X���LqE��9���;8C <���;�9LqE�X�����e��=��'��`c1�]�_�mF��;u��`   `   j�n�|g��0Q�A`1�{���RѽOя��1��ɷ�����];5<L
9<5<��];���ɷ��1�Oя��Rѽ{��A`1��0Q�|g�`   `   	3��;-����6/�@eӽ���S�K���|zf����P�;k9<؛R<k9<�P�;��|zf�K���S����@eӽ6/�����;-�`   `   %���!@��P�ݽ�ͻ�����zW�wk�F��?ͻ��D;V<'�S<�g<'�S<V<��D;?ͻF��wk�zW������ͻ�P�ݽ!@��`   `   ���]o��%p����s�GZ<�8��H򞼊G
�C�9���;�8<�b<�wo<�b<�8<���;B�9�G
�H�8��GZ<���s�%p��]o��`   `   �E�=,>��1)��)
��˼pC�����L"��1��;
<\�C<$F\<[�c<$F\<\�C<
<1��;N"�����pC���˼�)
��1)�=,>�`   `   �x���i���ؘ��>f���s�\�T)�:Xm�;�<��<ά0<
�8<�!;<
�8<ά0<��<�<Wm�;S)�:s�\����>f��ؘ��i��`   `    썻OIu��	��?�9�:;,��;�N�;L� <�<��;*,�;s��;(e�;s��;),�;��;�<L� <�N�;,��;�:;�?�9�	�OIu�`   `   �d<��<�<d�#<��)<��&<|k<� �;˩;��,;)۶9����~캙���%۶9��,;˩;� �;|k<��&<��)<d�#<�<��<`   `   ��<*�<�̉<���<9�j<�A<�<�|;"��[�ɻ��*�B�Y��j�B�Y���*�[�ɻ"���|;�<�A<9�j<���<�̉<*�<`   `   4b�<�0�<��<�<!�y<a�)<��;�[�	�;�
���l�ռ����w������l�ռ
���
�;��[���;a�)<!�y<�<��<�0�<`   `   D��<R=�<�X�<]\�<��\<@��;hS[�k��ּP���]C���^��8h���^��]C�Q���ּk�kS[�?��;��\<]\�<�X�<R=�<`   `   '�<�a�<pS�<	
�<�h<�Q{���e��\�a3<���~�M ��TW��75��TW��M ����~�a3<��\𼈸e��Q{��h<
�<pS�<�a�<`   `   ��<k��<~ܦ<l
^<H�_;t�)��{�O�E�G��T������9 �x���9 ���T���G��O�E��{�u�)�E�_;l
^<~ܦ<k��<`   `   j��<�}�<8�<�<�������5�~Y��>�ͽA%�;`�^\1���7�^\1�;`�A%�>�ͽY���5��������<8�<�}�<`   `   �a�<�z�<��^<��H;��P��E�:���=Ž3	��#0�?R�<�i��9r�<�i�?R��#0�3	��=Ž:���E���P���H;��^<�z�<`   `   V�<7D�<�<�B��뱼 |C�.��<U��1-�(�]��B���(��.����(���B��(�]�1-�<U��.�� |C��뱼�B��<7D�<`   `   ��<��Z<���;R��\\����v���˽cs���O�C؄�᭞��°��H���°�᭞�C؄���O�cs���˽��v�\\��S�����;��Z<`   `   G�Y<��*<���:�e��`�]P��:,�b0-���l������7���ʾ�Ѿ�ʾ�7��������l�b0-�:,�]P���`��e���:��*<`   `   �M4<"	<ź������w0��Π��o �� <�q��4C�� �ľ�U۾z���U۾ �ľ4C��q��� <��o ��Π�w0�����˺��!	<`   `   ��<���;��W��t��5<�&��y#��(B�C������1ʾ�~�����~�1ʾ����C���(B�y#�&��6<��t����W����;`   `   #w<���;���O}���<�as���"c>��O��CԤ�K�ľ�e۾0�㾗e۾K�ľCԤ��O��"c>��as���<�P}��������;`   `   Z�<���;�[o��w��b0��������_1�Np�ᅘ������ʾ�Ѿ�ʾ����ᅘ�Np�_1��������b0��w���[o����;`   `   ��< �;d	�aޅ�˧�����>ٽ���S�W���,����"Զ���,��W����S����>ٽ���̧�aޅ�h	� �;`   `   :C <���;e�9JqE�W�����e��=��'��`c1�]�_�mF��;u��Í��;u��mF��]�_�`c1�'���=����e�W���KqE�G�9���;`   `   N
9<5<��];���ɷ��1�Oя��Rѽ{��A`1��0Q�|g�j�n�|g��0Q�A`1�{���RѽOя��1��ɷ�����];5<`   `   ۛR<n9<Q�;��yzf�I���
S����@eӽ6/�����;-�	3��;-����6/�@eӽ���
S�J���zzf���Q�;m9<`   `   �g<)�S<V<ȏD;?ͻF��vk�yW������ͻ�O�ݽ!@��%���!@��O�ݽ�ͻ�����zW�wk�F��?ͻÏD;V<)�S<`   `   Q�%<f�<���;}ɺ��;�i�̼�-��E���	���s۽	S����z����	S��s۽�	���E���-�i�̼��;��ɺ���;f�<`   `   �<Q�<�%�;4; }��\�Q���ü��rS�T���[������ ��������[��U��rS�����ü]�Q�"}��
4;�%�;P�<`   `   ��;Ȓ�;�Í;'�/;�|H��H��a+.�!���h�ڼS����.�p�C�D�J�p�C���.�S��h�ڼ!���b+.��H���|H�$�/;�Í;Ȓ�;`   `   &�
����=��v ݹ�b���2�fl�~0���O�9�\��ƍ����z������ƍ�9�\��O��0��il��2�:c��� ݹ"=�����`   `   �bo�a�a�;�;���B���Lഺ2]h:r ;��:.o�:�%(��}��C���}�%&(�*o�:��:r ;&]h:RഺC�����;�;�a�a�`   `   `�
�A��0��T����j��
�hO7�P�;#.�;,� <��2<":<�;<":<��2<+� <".�;
P�;rO7��
维�j��T���0�A�`   `   U1}�>"s���V���,�L����є������:��<hub<��<���<�<���<��<hub<��<��:��뻨є�L�����,���V�>"s�`   `   ��νkVǽ�ᱽ|I����Z��|����c��t��;D/f<v��<p��<��<p��<v��<D/f<s��;c������|���Z�|I���ᱽkVǽ`   `   ���\M�+���"�.���u@q��t��k}��ᄷ��7<�՘<�N�<�k�<�N�<�՘<��7<+ℷ�k}��t�u@q�.����"�+��\M�`   `   �e� ]��{F�w�%�� ��ﶽc�h�Mq��ҵ��z�;�	�<�3�<�<�3�<�	�<�z�;ӵ�Mq��c�h��ﶽ� �w�%��{F� ]�`   `   �'��1���1ǉ��]f��J3�J�Q��ZC��!��<e��m0<<��<x�<��<m0<<<e���!��ZC�Q��J��J3��]f�1ǉ�1���`   `   QMԾ��̾@���ݘ���m��{,���潐Ί��
��z��n�;R�s<��<R�s<�n�;�z��
��Ί�����{,���m��ݘ�@����̾`   `   δ�D���O�<������?gZ��n���jFC�������7Ic,<t�c<Ic,<��7����jFC��𵽐n�?gZ����<����O�D��`   `   ��%��<���G��7l���y���;2�vM߽,�y�æ�'o»il�;ϲ"<il�;'o»æ�,�y�vM߽�;2��y��7l��G�����<�`   `   >�?�pd8��#����о�~���mL�$C��]��^=��8�;n�;;�8�^=��]��$C��mL��~��о����#�pd8�`   `   �NR�X�I��2��'�vX�������^�	��"W����'��J}�텯�ΊO;텯��J}���'�"W��	����^�����vX⾗'��2�X�I�`   `   ��X��'P�Ld8����N�9֨�Yf��e��䭽�5�9@����n�%x:��n�9@���5��䭽�e�Yf�9֨��N���Ld8��'P�`   `   KR��I��3�Y�����zB���Yb������N�6��I�������3�����I��N�6�������Yb�zB�����Y���3��I�`   `   ��?��d8�  $�״�jWҾ���QS���������,��R�����L����R����,�������QS����jWҾ״�  $��d8�`   `   �D%������lS�BX��>h���r;���t��z�ZN{�� J�?�^:� J�ZN{�z�t�����r;�>h��BX��lS쾪����`   `   �����Q�mcþ����-c�����ͽ�s�/��6;�.n<�)�2;.n<�6;�/���s��ͽ���-c�����mcþ�Q��`   `   ��ѾÚʾ{w��콙��0s�W�4�*C��~-��`=>�����޻�;H��;�;�޻���`=>�~-��*C��W�4��0s�콙�{w��Úʾ`   `   Q�������H
���df��7�t���0���/s����xFo��5�C@�;zu�;C@�;�5�xFo�����/s��0��t���7��df�H
������`   `   JB\��U�A�|�#�����S½����
'��ܯ�M5�\�;���;<���;\�;M5�ܯ��
'�����S½���|�#�A��U�`   `   z����
S��s۽�	���E���-�j�̼��;��ɺ���;c�<N�%<c�<���;�ɺ��;�j�̼�-��E���	���s۽
S����`   `    ��������[��U��rS�����ü_�Q�&}��4;�%�;N�<�<N�<�%�;4;&}��_�Q���ü��rS�U���[������`   `   E�J�q�C���.�T��i�ڼ"���d+.��H��_}H��/;�Í;Ē�;��;Ē�;�Í;�/;b}H��H��d+.�"���i�ڼT����.�q�C�`   `   z������ƍ�<�\��O��0��ql�2�(d��� ݹ1=��ǉ�.�
�ǉ�1=��� ݹ4d�� 2�rl��0���O�<�\��ƍ����`   `   �C���}��((�o�:Թ�:r ;]h:aഺG�����=�;�c�a��bo�c�a�=�;���G���bഺ]h:r ;ӹ�:o�:�((��}�`   `   �;<:<��2<)� <.�;P�;�O7��
绶�j��T���0�A�`�
�A��0��T����j��
绒O7�P�;.�;)� <��2<:<`   `   �<���<��<fub<��<��:��뻩є�M�����,���V�>"s�U1}�>"s���V���,�M����є������:��<fub<��<���<`   `   ��<o��<u��<B/f<p��;f������|���Z�|I���ᱽkVǽ��νkVǽ�ᱽ|I����Z��|����g��p��;B/f<u��<o��<`   `   �k�<�N�<�՘<��7<�䄷�k}��t�v@q�/����"�+��\M����\M�+���"�/���v@q��t��k}��儷��7<�՘<�N�<`   `   �<�3�<�	�<�z�;ӵ�Nq��c�h��ﶽ� �w�%��{F� ]��e� ]��{F�w�%�� ��ﶽc�h�Nq��Ե��z�;�	�<�3�<`   `   x�<��<m0<<Be���!��ZC�Q��J��J3��]f�1ǉ�1����'��1���1ǉ��]f��J3�J�Q���ZC��!��Fe��l0<<��<`   `   ��<R�s<�n�;�z��
��Ί�����{,���m��ݘ�@����̾QMԾ��̾@���ݘ���m��{,���潐Ί��
��z��n�;R�s<`   `   t�c<Ic,<��7����kFC��𵽐n�@gZ����<����O�D��δ�D���O�<������@gZ��n���kFC�������7Ic,<`   `   ϲ"<il�;&o»¦�,�y�vM߽�;2��y��7l��G�����<���%��<���G��7l���y���;2�vM߽-�y�æ�'o»il�;`   `   n�;;�8�^=��]��$C��mL��~��о����#�pd8�>�?�pd8��#����о�~���mL�$C��]��^=��8�;`   `   ҊO;兯��J}���'�"W��	����^�����vX⾘'��2�X�I��NR�X�I��2��'�vX�������^�	��"W����'��J}�煯�`   `   9x:��n�8@���5��䭽�e�Yf�9֨��N���Ld8��'P���X��'P�Ld8����N�9֨�Yf��e��䭽�5�9@����n�`   `   ��3�����I��N�6�������Yb�zB�����Y���3��I�KR��I��3�Y�����zB���Yb������N�6��I�����`   `   ��L����R����,�������QS����jWҾ״�  $��d8���?��d8�  $�״�jWҾ���QS���������,��R����`   `   `�^:� J�XN{�z�t�����r;�>h��BX��lS쾪�����D%������lS�BX��>h���r;���t��z�YN{�� J�`   `   2�2;n<�4;�/���s��ͽ���-c�����mcþ�Q�������Q�mcþ����-c�����ͽ�s�/��5;�n<�`   `   L��;�;�޻���_=>�~-��)C��W�4��0s�콙�{w��Úʾ��ѾÚʾ{w��콙��0s�W�4�*C��~-��_=>�����޻�;`   `   u�;H@�;�5�uFo�����/s��0��t���7��df�H
������Q�������H
���df��7�t���0���/s����vFo��5�G@�;`   `   <���;g�;G5�ܯ��
'�����S½���|�#�A��U�JB\��U�A�|�#�����S½����
'��ܯ�I5�d�;���;`   `   ��;�+L;8����?�`+ռ��;��}����ѽ�?���/�2�N�0yd��'l�0yd�2�N���/��?���ѽ�}����;�`+ռ��?�;���+L;`   `   c)\;��;�!_��ڻ���Q�^�6�����8���^޽1���&�G���&�1���^޽�8�����_�6�Q缮���ڻ�!_���;`   `   8\��?=�vp^�7���{�$�Ġ���Ѽ�,���K�g����ϗ�����:P�������ϗ�h�����K��,��ѼŠ��|�$�8���xp^�A=�`   `   ܪL�J�F�.�7�R�(�ϣ$��Z6�cd����}&ɼÃ��R`��7(��C.��7(�R`�Ã��}&ɼ���cd��Z6�У$�R�(�/�7�J�F�`   `   �n����#ռǪ��䔇���I�.��#�u��)�L8I�!�b�� l�!�b�L8I�)�v��#�/����I�䔇�Ǫ��#ռ��`   `   ̣o�X�f�?M�MC(�����h⨼*C��p���*O����:F;~�b;�Nh;}�b;F;���:�*O��p��+C�i⨼����MC(�?M�X�f�`   `   y`ͽe�Ž���u��^����l������s;:���;Ԫ9<]<0�g<]<Ԫ9<���;�s;:����l����^��u����e�Ž`   `   �<$��p��*�W���� �~����m����Z�c�;O�k<ߖ�<���<ߖ�<O�k<c�;��Z�m����� �~���W���*��p�`   `   �4z�*_q��X�V�4�;�Ƚm���N����H�2�Y;R]<�=�<�,�<�=�<R]<2�Y;��H�N��m���Ƚ;�V�4��X�*_q�`   `   �L��x����W������!M�y����½�-c��Rмyo��u�<��<^�<��<u�<yo���Rм�-c���½y���!M�����W��x���`   `   �������޾I��JR����N�5a
�K�����,��lk�X�i;�]<A��<�]<X�i;�lk���,�K���5a
���N�JR��I����޾���`   `   -�0�)�)�@��{��_��������9�Ί��q{�ؼ����
<��J<
<����ؼ�q{�Ί彶�9����_���{��@��)�)�`   `   Khg�Z�]�"D��� �C������ol�w��Ì��S� ��	H��+;��;�+;�	H�S� �Ì��w��ol�����C���� �"D�Z�]�`   `   d����[��`s�cnE�y��M�Ծ�Ǝ���3�н:T�5+���3W��6;�3W�5+��:T�н��3��Ǝ�M�Ծy��cnE�`s��[��`   `   ���_��cŎ��Pf�B-�A��#���N���w��.�	X��/�	X�.㼶w�����N�#��A��B-��Pf�cŎ�_��`   `   ���<��g֝��t}���=����0貾�Db�M�T"��@��Y�U�h�ػY�U�@��T"��M��Db�0貾�����=��t}�g֝�<��`   `   M�ĿdŻ��^��k���D�>K
�E
��U�j��,�J(��K������6������K��J(���,�U�j�E
��>K
��D�k���^��dŻ�`   `   g���D������~���>��
��s��tg�X�����EI����-���EI�����X�tg��s���
���>��~�����D��`   `   g����^�����Egg��.��|���Ũ���X�y��pW�����熼W�(��熼��pW��y����X��Ũ��|���.�Egg�����^��`   `   U��g6���ps�2�F����hھ�
��ɪ@����市��C��`h� ���`h��C�市����ɪ@��
���hھ��2�F��ps�g6��`   `   Qf��]��D���!��~��ݞ���2z���"�l�Ž]�[���Լe�.�����e�.���Լ]�[�l�Ž��"��2z�ݞ���~����!��D��]�`   `   -�.�@Z(��Q�p?���[þ����z�G�E{�v%��=,�qL��5�һ�5�һqL��=,�v%��E{�z�G������[þp?���Q�@Z(�`   `   TM��^E���Zܾ���\ꑾ�X��x�,�Ž�Um�=R��սJ������:���սJ�=R���Um�,�Ž�x��X�\ꑾ����Zܾ^E��`   `   �6���:������xĂ���O�e5��jٽ�>���%�������ѻ�B�:bu;�B�:��ѻ�����%��>���jٽe5���O�xĂ������:��`   `   �'l�1yd�3�N���/��?���ѽ�}����;�a+ռ��?�C���+L; ��;�+L;C����?�a+ռ��;��}����ѽ�?���/�3�N�1yd�`   `   G���&�1���^޽�8�����_�6�Q缰���ڻ�!_���;Z)\;��;�!_��ڻ���Q�_�6�����8���^޽1���&�`   `   :P�������ϗ�h�����K��,��ѼƠ��~�$�<����p^�H=�H\��H=��p^�<���~�$�Ơ���Ѽ�,���K�h����ϗ�����`   `   �C.��7(�R`�Ń��~&ɼ���cd��Z6�ң$�T�(�1�7�L�F�ުL�L�F�1�7�T�(�ң$��Z6�cd����~&ɼŃ��R`��7(�`   `   � l�#�b�N8I�Ō)�x��	#�1����I�唇�Ȫ��#ռ���n����#ռȪ��唇���I�1��	#�x��Ō)�N8I�#�b�`   `   �Nh;t�b;F;��:�*O��p��-C�j⨼����MC(�?M�Y�f�ͣo�Y�f�?M�MC(�����j⨼-C��p���*O���:F;s�b;`   `   .�g<]<Ҫ9<}��;�s;:����l����^��u����e�Žz`ͽe�Ž���u��^����l������s;:}��;Ҫ9<]<`   `   ���<ޖ�<M�k<_�;��Z�m����� �~���X���*��p��<$��p��*�X���� �~����m����Z�_�;M�k<ޖ�<`   `   �,�<�=�<R]<,�Y;��H�N��m���Ƚ;�V�4��X�*_q��4z�*_q��X�V�4�;�Ƚm���N����H�+�Y;R]<�=�<`   `   ^�<��<t�<|o���Rм�-c���½y���!M�����W��x����L��x����W������!M�y����½�-c��Rм|o��s�<��<`   `   @��<�]<U�i;�lk���,�K���5a
���N�JR��I����޾����������޾I��JR����N�5a
�K�����,��lk�T�i;�]<`   `   ��J<
<����ؼ�q{�Ί彷�9����_���{��@��)�)�-�0�)�)�@��{��_��������9�Ί��q{�ؼ����
<`   `   ��;�+;�	H�S� �Ì��w��ol�����C���� �"D�Z�]�Khg�Z�]�"D��� �C������ol�w��Ì��T� ��	H��+;`   `   �6;�3W�4+��:T�н��3��Ǝ�M�Ծy��cnE�`s��[��d����[��`s�cnE�y��M�Ծ�Ǝ���3�н:T�5+���3W�`   `   �/�X�.㼵w�����N�#��A��B-��Pf�cŎ�_�����_��cŎ��Pf�B-�A��#���N���w��.�X�`   `   f�ػX�U�@��T"��M��Db�0貾�����=��t}�g֝�<�����<��g֝��t}���=����0貾�Db�M�T"��@��X�U�`   `   5������J��J(���,�U�j�E
��>K
��D�k���^��dŻ�M�ĿdŻ��^��k���D�>K
�E
��U�j��,�J(��J������`   `   �-���DI�����X�tg��s���
���>��~�����D��g���D������~���>��
��s��tg�X�����EI���`   `   U�(��熼��pW��y����X��Ũ��|���.�Egg�����^��g����^�����Egg��.��|���Ũ���X�y��pW�����熼`   `   ���`h��C�市����ɪ@��
���hھ��2�F��ps�g6��U��g6���ps�2�F����hھ�
��ɪ@����市��C��`h�`   `   ����c�.���Լ]�[�l�Ž��"��2z�ݞ���~����!��D��]�Qf��]��D���!��~��ݞ���2z���"�l�Ž]�[���Լc�.�`   `   �0�һpL��=,�v%��E{�z�G������[þp?���Q�@Z(�-�.�@Z(��Q�p?���[þ����z�G�E{�v%��=,�pL��1�һ`   `   �:���ҽJ�;R���Um�+�Ž�x��X�\ꑾ����Zܾ^E��TM��^E���Zܾ���\ꑾ�X��x�+�Ž�Um�<R��ӽJ����`   `   ku;C�:��ѻ�����%��>���jٽe5���O�xĂ������:���6���:������xĂ���O�e5��jٽ�>���%�������ѻ�B�:`   `   ��h�!�P�s�)��½�I1/����~ڽ���D�N�'������ ��1��� �����'��D�N�����~ڽ��I1/��½�t�)�"�P�`   `   �	;��f�����Y�������<�e���;�ǽ�^�5`%��JB�.>V��a]�.>V��JB�5`%��^�;�ǽf�����<�����Y�����f��`   `   e"��)��3D�G{�六��(���;0��Fr���qŽ%"�}P���K�}P��%"�qŽ�𞽼Fr��;0��(��六�H{��3D��)�`   `   �Ƽ�!¼&���녯�t����6��3,������/���V���y��L��߸���L����y���V���/����3,༘6��u���셯�&����!¼`   `   �~G��A��2/��K�$��(�˼'3��e5���/���ȼ�G������]�������Gἐȼ�/��f5��'3��(�˼$���K��2/��A�`   `   ����i�����%Ȃ��zL��i�i�ͼو�ƨ8����="뻛�ỂaỜ��="뻃��ƨ8�و�j�ͼ�i��zL�%Ȃ�����i��`   `   ����a����7|ڽ�s��;Ar�a1�<'��Q�����nm;���;q��;���;�nm;����Q�<'��a1�;Ar��s��7|ڽ����a�`   `   ;�p�-h�eoP�m5.�E�+½YX}��9�۵y�M��H6�;��I<�tb<��I<G6�;M��۵y��9�YX}�+½E�m5.�eoP�-h�`   `   m)���w��⟾G����N�,�lŽ%@i��(ἇ�㻡r�;�o\<u�<�o\<�r�;����(�%@i�lŽ,���N�G��⟾�w��`   `   �3
�����1��ľWݗ��Z��'�Ӽ���:��狼�m�:G�5<C�i<G�5<�m�:�狼�:�Ӽ���'��Z�Wݗ���ľ�1����`   `   +VH�P@��j*����{־R�����M�D��h�������߻Ab�;y*<Ab�;�߻���h���D����M�R����{־���j*�P@�`   `   ������:�l�QT@�K����ξ�Љ�՟+��rý�a@��r��E�f��;E�f��r���a@��rý՟+��Љ���ξK��QT@�:�l����`   `   �f��Ù��)����}��h=�����	����[�%5��.ރ�ѭ�N����|��N���ѭ�.ރ�%5����[��	������h=���}�)��Ù��`   `   ���N���ɿ�v��K�j���"��־"H������Ȧ���f�t�����f�t����Ȧ����"H���־��"�K�j��v���ɿN��`   `   ���}���򿬞������Fg=��:��H���ȕ4��DŽ��B��W��ީ]��W����B��DŽȕ4�H����:��Fg=�����������}��`   `   �*��� �V��iӿ����]P��E�{��VfF�^�۽��`�J
ݼ7���J
ݼ��`�^�۽VfF�{���E�]P������iӿV��� �`   `   Ԧ1�$�'�$����ۿ8��S]W����C����N��f罅�q�����I�������q��f罝�N��C����S]W�8����ۿ$��$�'�`   `   S*�8� ��s���ӿ5?���Q�����^����L����ԣt��� �J5���� �ԣt���潢�L��^������Q�5?����ӿ�s�8� �`   `   �����7���e��_&���M@������۟�H9@�Vڽ0�h�&_���²�&_��0�h�VڽH9@��۟������M@�_&���e��7����`   `   !���Ў�v�ɿW����m���&�J޾	�����+��ý"�P�=�ۼr��=�ۼ"�P��ý��+�	���J޾��&���m�W��v�ɿЎ�`   `   j������v��J��N@�y��f&��Hcn�SX��ץ���.������y������.��ץ�SX�Hcn�f&��y���N@�J�v�����`   `   At������p�k�A*A��
�8־�ђ�
�>��������"��蘃�-�蘃�"���������
�>��ђ�8־�
�A*A�p�k�����`   `   F�D��h=�x�(�N���پ�៾�]��_�C��riG���ļ1)�%û1)���ļriG�C���_��]��៾��پN�x�(��h=�`   `   � ��U��=���¾O���d�0���2ҽ�/����|����T�����T��|������/���2ҽ0��d�O�����¾�=辂U�`   `   1��� �����'��D�N�����~ڽ��J1/��½�v�)�*�P��h�*�P�v�)��½�J1/����~ڽ���D�N�'������ ��`   `   �a]�.>V��JB�5`%��^�<�ǽf�����<�����Y�����f���	;��f�����Y�������<�f���<�ǽ�^�5`%��JB�.>V�`   `   �K�~P��%"�qŽ�𞽽Fr��;0��(��慭�J{��3D��)�g"��)��3D�I{�慭��(���;0��Fr���qŽ%"�~P��`   `   ߸���L����y���V���/����4,༙6��v���텯�'����!¼�Ƽ�!¼'���텯�v����6��4,������/���V���y��L��`   `   �]�������Gἑȼ�/��g5��(3��)�˼$���K��2/��A��~G��A��2/��K�$��)�˼(3��g5���/���ȼ�G�����`   `   �aỠ��B"뻅��Ȩ8�و�k�ͼ�i��zL�%Ȃ�����i������i�����%Ȃ��zL��i�k�ͼو�Ȩ8����B"뻠��`   `   m��;���;�nm;����Q�='��a1�;Ar��s��7|ڽ����a�����a����7|ڽ�s��;Ar�a1�='��	Q������nm;���;`   `   �tb<��I<D6�;'M��ݵy��9�YX}�,½E�m5.�foP�-h�;�p�-h�foP�m5.�E�,½YX}��9�ݵy�(M��C6�;��I<`   `   t�<�o\<�r�;����(�%@i�lŽ,���N�G��⟾�w��m)���w��⟾G����N�,�lŽ%@i��(Ἂ�㻝r�;�o\<`   `   A�i<F�5<�m�:�狼�:�Ӽ���'��Z�Wݗ���ľ�1�����3
�����1��ľWݗ��Z��'�Ӽ���:��狼�m�:F�5<`   `   x*<@b�;�߻���h���D����M�R����{־���j*�P@�+VH�P@��j*����{־R�����M�D��h�������߻?b�;`   `   췢;e�f��r���a@��rý՟+��Љ���ξL��RT@�:�l����������:�l�QT@�L����ξ�Љ�՟+��rý�a@��r��l�f�`   `   �|��O���ҭ�.ރ�%5����[��	������h=���}�)��Ù���f��Ù��)����}��h=�����	����[�%5��.ރ�ҭ�O���`   `   ����f�t����Ȧ����"H���־��"�K�j��v���ɿN�����N���ɿ�v��K�j���"��־"H������Ȧ���f�t�`   `   ީ]��W����B��DŽȕ4�H����:��Fg=�����������}�����}���򿬞������Fg=��:��H���ȕ4��DŽ��B��W��`   `   6���J
ݼ��`�^�۽VfF�{���E�]P������iӿV��� ��*��� �V��iӿ����]P��E�{��VfF�^�۽��`�J
ݼ`   `   �I�������q��f罝�N��C����S]W�8����ۿ$��$�'�Ԧ1�$�'�$����ۿ8��S]W����C����N��f罅�q����`   `   I5���� �ԣt���潢�L��^������Q�5?����ӿ�s�8� �S*�8� ��s���ӿ5?���Q�����^����L����ԣt��� �`   `   �²�%_��0�h�VڽH9@��۟������M@�_&���e��7���������7���e��_&���M@������۟�H9@�Vڽ0�h�%_��`   `   r��<�ۼ!�P��ý��+�	���J޾��&���m�W��v�ɿЎ�!���Ў�v�ɿW����m���&�J޾	�����+��ý!�P�<�ۼ`   `   ��y������.��ץ�SX�Hcn�f&��y���N@�J�v�����j������v��J��N@�y��f&��Hcn�SX��ץ���.����`   `   -�瘃�!���������	�>��ђ�8־�
�A*A�p�k�����At������p�k�A*A��
�8־�ђ�	�>��������"��瘃�`   `    û1)���ļqiG�C���_��]��៾��پN�x�(��h=�F�D��h=�x�(�N���پ�៾�]��_�C��qiG���ļ1)�`   `   ���T��z������/���2ҽ0��d�O�����¾�=辂U�� ��U��=���¾O���d�0���2ҽ�/����{����T��`   `   Ҹֻ�$��_��$��ax�>�ƽ�A���S��������e�վ��wV����e�վ���������S��A�>�ƽax�%���_���$�`   `   �-�,�0�u���қؼ��-�{݅�d�Ľ��	��#6���c�;0��F��:V��F��;0����c��#6���	�d�Ľ{݅���-�ӛؼu���,�0�`   `    f��#q���ܩ�*μr��$�8�ez~�N֫�3<߽��	��/!�e>1�W�6�e>1��/!���	�3<߽N֫�ez~�$�8�s��*μ�ܩ�$q��`   `   ����?�y������4�Б�'�,���S��т���������ǽ�5ͽ�ǽ��������т���S�'�,�Б��4����y���?�`   `   ez��XV���x���X�/�8��R��H�k`�&�0j(��J;�F�I��O�F�I��J;�0j(�&�l`��H��R�/�8���X��x�XV��`   `   N������ֽ�u������]���#�����#ļ�Q��z�����G,�����z���Q��#ļ������#��]�����u���ֽ��`   `   >yL�fE�f�1��B�vC�1׫�I�k��&��t���M�V�ш��[�ш�V��M��t���&�I�k�2׫�vC��B�f�1�fE�`   `   G���֪���R����m�+X9�����r���_����}VS�Q����O;��;��O;R��}VS�����_��r�����+X9���m��R��֪��`   `   b� �����4ݾ������J;M�1�	�0����B;�I��!i���F�;�}�;�F�;!i��I���B;�0���1�	�J;M��������4ݾ���`   `   s�D���<�8['�,�	��Ҿ�ꖾJJ�̟���ʍ�{����,��G�:s��;�G�:��,�{���ʍ�̟��JJ��ꖾ�Ҿ,�	�8['���<�`   `   �ᒿ����o�v���G����i�վ�5��M;1���˽,�N�u���*r��v�v:*r��v���,�N���˽M;1��5��i�վ�����G�o�v�����`   `   n�տ�˿>����ˌ���P��w�|u����m��
�+ܑ�s����@��4����@�s��+ܑ��
���m�|u���w���P��ˌ�>����˿`   `   y�����@���׾������=��T���	���21�%���n ;�0Ħ���L�0Ħ�n ;�%����21��	���T����=�����׾��@����`   `   �XL�,<@�_i!�p���gk��O�k�������W����L�p��������L�p������W�����O�k�gk��p���_i!�,<@�`   `   �c����s���H��s�ٸѿ)����/�Z�վ�)y��	�*��ζ��[ؼζ�)���	��)y�Z�վ�/�)���ٸѿ�s���H���s�`   `   sc��am���g�S�*��꿁|����@���;���	0�t顽Ru/�ؗ�Ru/�t顽	0�;����꾙�@��|����S�*��g�am��`   `   �}�� ����s��x2�\?��Z=����G�X������G������">�����">������G����X���G�Z=��\?���x2��s� ���`   `   �a���q����g�>+����ֈ���#C�B�����5���VA��P�VA����5����B��#C�ֈ�����>+���g��q��`   `   �W���s�K7I�����Nӿ䁌��3��,ݾ�5���,��)��=8����=8��)���,��5���,ݾ�3�䁌��Nӿ���K7I��s�`   `   �L�a@�Η!�r����X��bnp� �v�¾�hi�����T��A�$�K��A�$��T������hi�v�¾ �bnp��X��r���Η!�a@�`   `   �s����?���ӿ�������B�� ��
���YE�}����w��\	��nͼ�\	���w�}���YE��
��� ���B������ӿ��?����`   `   A@ԿE]ʿ���W��a�S���2ʾ[ꁾȱ�|���2jE�E�Լ�1��E�Լ2jE�|���ȱ�[ꁾ2ʾ��a�S�W�����E]ʿ`   `   _���}���U�t�c�G�� 3ݾ�����aE�����l�����X'���U�X'������l������aE����� 3ݾ�c�G�U�t�}���`   `   6�?��88�xB$� u���ԾoH���tY����밽��J���ҼΎN�c�	�ΎN���Ҽ��J��밽���tY�oH����Ծ u�xB$��88�`   `   wV����e�վ���������S��A�>�ƽax�%���_���$�ָֻ�$��_��%��ax�>�ƽ�A���S��������e�վ��`   `   :V��F��;0����c��#6���	�d�Ľ{݅���-�ԛؼv���.�0��-�.�0�v���ԛؼ��-�{݅�d�Ľ��	��#6���c�;0��F��`   `   W�6�e>1��/!���	�4<߽N֫�fz~�%�8�s��+μ�ܩ�$q��!f��$q���ܩ�+μs��%�8�fz~�N֫�4<߽��	��/!�e>1�`   `   �5ͽ�ǽ��������т���S�(�,�Б��4����y���?�����?�y������4�Б�(�,���S��т���������ǽ`   `   �O�F�I��J;�1j(�&�l`��H��R�/�8���X��x�XV��ez��XV���x���X�/�8��R��H�l`�&�1j(��J;�F�I�`   `   H,�����z���Q��$ļ������#��]�����u���ֽ��N������ֽ�u������]���#�����$ļ�Q��z�����`   `   �[�ш��V��M��t���&�I�k�2׫�wC��B�f�1�fE�>yL�fE�f�1��B�wC�2׫�I�k��&��t���M��V�ш�`   `   ��;��O;Y��VS�����_��r�����+X9���m��R��֪��G���֪���R����m�+X9�����r���_����VS�Y����O;`   `   �}�;�F�;$i��I���B;�0���1�	�J;M��������4ݾ���b� �����4ݾ������J;M�1�	�0����B;�I��$i���F�;`   `   p��;�G�:��,�{���ʍ�̟��JJ��ꖾ�Ҿ,�	�8['���<�s�D���<�8['�,�	��Ҿ�ꖾJJ�̟���ʍ�{����,��G�:`   `   h�v:,r��v���,�N���˽M;1��5��i�վ�����G�o�v������ᒿ����o�v���G����i�վ�5��M;1���˽,�N�v���,r��`   `   �4����@�s��,ܑ��
���m�}u���w���P��ˌ�>����˿n�տ�˿>����ˌ���P��w�|u����m��
�,ܑ�s����@�`   `   ��L�1Ħ�n ;�%����21��	���T����=�����׾��@����y�����@���׾������=��T���	���21�%���n ;�1Ħ�`   `   �����L�p������W�����O�k�gk��p���_i!�,<@��XL�,<@�_i!�p���gk��O�k�������W����L�p���`   `   �[ؼζ�)���	��)y�Z�վ�/�)���ٸѿ�s���H���s��c����s���H��s�ٸѿ)����/�Z�վ�)y��	�)��ζ�`   `   ؗ�Ru/�t顽	0�;����꾙�@��|����S�*��g�am��sc��am���g�S�*��꿁|����@���;���	0�t顽Ru/�`   `   ����">������G����X���G�Z=��\?���x2��s� ����}�� ����s��x2�\?��Z=����G�X������G������">�`   `   �P�UA����5����B��#C�ֈ�����>+���g��q���a���q����g�>+����ֈ���#C�B�����5���UA�`   `   ���=8��)���,��5���,ݾ�3�䁌��Nӿ���K7I��s��W���s�K7I�����Nӿ䁌��3��,ݾ�5���,��)��=8�`   `   J��@�$��T������hi�v�¾ �bnp��X��r���Η!�a@��L�a@�Η!�r����X��anp� �v�¾�hi�����T��@�$�`   `   �nͼ�\	���w�}���YE��
��� ���B������ӿ��?�����s����?���ӿ�������B�� ��
���YE�}����w��\	�`   `   �1��D�Լ1jE�|���ȱ�[ꁾ2ʾ��a�S�W�����E]ʿA@ԿE]ʿ���W��a�S���2ʾ[ꁾȱ�|���1jE�D�Լ`   `   �U�W'������l������aE����� 3ݾ�c�G�U�t�}���_���}���U�t�c�G�� 3ݾ�����aE�����l�����W'��`   `   a�	�̎N���Ҽ��J��밽���tY�oH����Ծ u�xB$��88�6�?��88�xB$� u���ԾoH���tY����밽��J���Ҽ̎N�`   `   �3>�:�w�CeּC�=��8��R���S�=��-��񕶾���[�&��	�!�&���[���񕶾�-��S�=�R����8��C�=�Ceּ:�w�`   `   |Co����c?���*�d�e鬽P����70�_�i�[ƒ��y���.��T�ƾ�.���y��[ƒ�_�i��70�P���e鬽d��*�c?�����`   `    
м�yּ�켘j���5�{/u��9��[��?�*Y3���Q�+�f�n�+�f���Q�*Y3��?�[��9��{/u���5��j��켑yּ`   `   �C�k@�Z:��5�R�8���I��Rl��J��;,���}Խwd��u\��`	�u\�wd���}Խ;,���J���Rl���I�R�8��5�Z:�k@�`   `   ʍ�������<�������0u���X�\�J��?M��^���w��G��P�����P���G����w��^��?M�]�J���X��0u������<������`   `   s��h��ۥ�w���A������<f�~�9�~� ��F�N9�u@����u@�N9��F�~� �~�9��<f�����A��w��ۥ�h��`   `   �t����y�o+a��=���*_ཱི ��M^�Xb�f�༢H��k����m��l����H��f��Xb�N^�� ��*_ཪ��=�o+a���y�`   `    �Ҿ;˾t⵾�ȗ��l���-����W`��zB�3�缰뉼�h2�����h2��뉼4��zB�W`�������-��l��ȗ�t⵾;˾`   `   V�'�Ac!��|�_��(�������\3��G��G��R���������m!ֻ�������R���G���G��\3����(���_���|�Ac!�`   `   :y��1�{�m�]��4�r��Z�¾ł�1o%�6mĽ7]X���ټ��P�+7
���P���ټ7]X�6mĽ1o%�ł�Z�¾r���4�m�]�1�{�`   `   $�ʿ�2���ا��&���G�]������f��X�����B�G��:�X�G���B�����X���f����]��G��&���ا��2��`   `   ���U�����O���\���5%@�N���*��0k5���ɽ�"T�KX�l���KX��"T���ɽ0k5��*��N��5%@�\���O������U��`   `   \�d���V���2�X��m㾿0~��!��6ž��f�<� �y%��L1�� �L1�y%��<� ���f��6ž�!�0~�m㾿X����2���V�`   `   ?���_����w�e'5����L7����G���E���b���Ч��<�����<��Ч�b��E�������G�L7�����e'5���w�_��`   `   ����ɟ���G��d�a��>⾿�j�=Y�aˠ�aE3���½��]��V*���]���½aE3�aˠ�=Y��j�>⾿a��d��G��ɟ��`   `   e�&� ��6������+�+.տjI�����j믾�LD��YֽR�v��?�R�v��Yֽ�LD�j믾���jI��+.տ�+�����6��&� �`   `   H��s�
���������2�%�ݿ$����������>L�!�R�&=J�R�!ཪ>L��������$��%�ݿ�2��������s�
�`   `   �c�*� ��Q���ӄ�9�+��wֿ.���'�������I��޽룁�=J�룁��޽��I�����'�.����wֿ9�+��ӄ��Q��*� �`   `   ��������to��Z�d�v���0��ױn�Ax�=�����=���ѽ3�t�~�>�3�t���ѽ��=�=���Ax�ױn��0��v��Z�d�to������`   `   Xx��\F��(x�7�5��k�������M�3���f���.)���1Z�^�)��1Z���.)��f��3����M�����k��7�5�(x�\F��`   `   �d�^V�T�2�'��1�������'���о��y�jy� ��*7��*7� ��jy���y���о��'�����1��'�T�2�^V�`   `   ���3�������¿�����hE��~��N���`H��P��E��Q��ۼ�Q��E��P罙`H��N���~��hE������¿����3��`   `   �ȿ�⾿R����%��9�I�S{�������y�9��~��A9B�S+ּ3*��S+ּA9B��~��9���y�����S{�9�I��%��R����⾿`   `   l���hv��Z�M3��
���Ⱦh<��a�4��U�p����q��Ϛ��c��Ϛ��q�p����U�a�4�h<����Ⱦ�
�M3��Z��hv�`   `   	�!�&���[���񕶾�-��S�=�R����8��D�=�Deּ<�w��3>�<�w�DeּC�=��8��R���S�=��-��񕶾���[�&��`   `   T�ƾ�.���y��[ƒ�_�i��70�P���f鬽d��*�d?�����}Co����d?���*�d�f鬽P����70�_�i�[ƒ��y���.��`   `   n�+�f���Q�*Y3��?�[��9��|/u���5��j�	�켒yּ 
м�yּ	�켘j���5�|/u��9��[��?�*Y3���Q�+�f�`   `   �`	�u\�xd���}Խ;,���J���Rl���I�S�8��5�Z:�k@��C�k@�Z:��5�S�8���I��Rl��J��;,���}Խxd��u\�`   `   ���P���G����w��^��?M�]�J���X��0u������<������ʍ�������<�������0u���X�]�J��?M��^���w��G��P��`   `   ���v@�O9��F�� ��9��<f�����A��w��ܥ�h��s��h��ܥ�w���A������<f��9�� ��F�O9�v@�`   `   �m��m����H��g��Yb�N^�� ��+_ཪ��=�o+a���y��t����y�o+a��=���*_ུ ��N^�Yb�g�༣H��m���`   `   ����h2��뉼4��zB�W`�������-��l��ȗ�t⵾;˾ �Ҿ;˾t⵾�ȗ��l���-����W`��zB�4�缱뉼�h2�`   `   p!ֻ�������S���G���G��\3�����(���`���|�Ac!�V�'�Ac!��|�`��(��������\3��G��G��S���������`   `   ,7
���P���ټ7]X�6mĽ1o%�ł�Z�¾r���4�m�]�1�{�:y��1�{�m�]��4�r��Z�¾ł�1o%�6mĽ7]X���ټ��P�`   `   ;�X�G���B�����X���f����]��G��&���ا��2��$�ʿ�2���ا��&���G�]������f��X�����B�G��`   `   l���KX��"T���ɽ0k5��*��N��5%@�\���O������U�����U�����O���\���5%@�N���*��0k5���ɽ�"T�KX�`   `   � �L1�z%��<� ���f��6ž�!�0~�m㾿Y����2���V�\�d���V���2�X��m㾿0~��!��6ž��f�<� �z%��L1�`   `   ����<��Ч�b��E�������G�L7�����e'5���w�_��?���_����w�e'5����L7����G���E���b���Ч��<�`   `   �V*���]���½aE3�aˠ�=Y��j�>⾿a��d��G��ɟ������ɟ���G��d�a��>⾿�j�=Y�aˠ�aE3���½��]�`   `   �?�R�v��Yֽ�LD�j믾���jI��+.տ�+�����6��&� �e�&� ��6������+�+.տjI�����j믾�LD��YֽR�v�`   `   &=J�R�!ཪ>L��������$��%�ݿ�2��������s�
�H��s�
���������2�%�ݿ$����������>L�!�R�`   `   =J�룁��޽��I�����'�.����wֿ9�+��ӄ��Q��*� ��c�*� ��Q���ӄ�9�+��wֿ.���'�������I��޽룁�`   `   }�>�3�t���ѽ��=�=���Ax�ױn��0��v��Z�d�to��������������to��Z�d�v���0��ױn�Ax�=�����=���ѽ3�t�`   `   ]�)��1Z���.)��f��3����M�����k��7�5�(x�\F��Xx��\F��(x�7�5��k�������M�3���f���.)���1Z�`   `   �*7����jy���y���о��'�����1��'�T�2�^V��d�^V�T�2�'��1�������'���о��y�jy����*7�`   `   �ۼ�Q��E��P罙`H��N���~��hE������¿����3�����3�������¿�����hE��~��N���`H��P��E��Q�`   `   2*��R+ּ@9B��~��9���y�����S{�9�I��%��R����⾿�ȿ�⾿R����%��9�I�S{�������y�9��~��@9B�R+ּ`   `   �c��Ϛ��q�p����U�a�4�h<����Ⱦ�
�M3��Z��hv�l���hv��Z�M3��
���Ⱦh<��a�4��U�p����q��Ϛ�`   `   ��~�����/���+d�����o��L�a�������۾1�j�)��>�&,F��>�j�)�1���۾����L�a�o�������+d�/������`   `   ׍��g���@��ۢ4��/���н��8�S��֌��^��SGҾ�v�O��v�SGҾ�^���֌�8�S����н�/��ۢ4�@��g���`   `   �j �q����I]/��*a��1���wͽ�t	���1�(Q[�[&��s��V���s��[&��(Q[���1��t	��wͽ�1���*a�I]/���q��`   `   �&i���f���a�x_�(�f��_�����P"��Ғὰ�����?�(�q�-�?�(�������Ғ�P"�������_�(�f�x_���a���f�`   `   yoѽ<̽Ɨ��!'��	3��.ŉ��-��Kb�����P��mY���ɽ�ν�ɽmY��P�����Kb���-��.ŉ�
3��!'��Ɨ��<̽`   `   6�5��=0�*� ��Q
��_佇���z���Z)���>n��Vk���q��y��M|��y���q��Vk��>n�Z)��z��������_佡Q
�*� ��=0�`   `   >G��o�����4�a��84��w	��&̽䗽z#k�M�C�Z)0�)c(�z&�)c(�Z)0�M�C�z#k�䗽�&̽�w	��84�4�a����o��`   `   ke�����tپ>d��R��0R�����Tͽg�����J�z��X�����X��z����J�g����Tͽ����0R�R�>d���tپ��`   `   �gL�e6D�$�-�����۾S5��BW[��Q��]��[�u��](��� �'�鼑� ��](�[�u��]���Q�BW[�S5����۾��$�-�e6D�`   `   i����_��!݈�Z]�m&���뾘ʞ�q�L�wD ������I�_��x���_���I�����wD �q�L��ʞ����m&�Z]�!݈��_��`   `   �������dԿ1�����u�w�)�ww߾���/K,�A�ν�^{��A(�4���A(��^{�A�ν/K,����ww߾w�)���u�1���dԿ����`   `   �jM�/JA��_"�$J���d��/�l���1���q�`�������FI�p�'�FI�������q�`�1�����/�l��d��$J���_"�/JA�`   `   as�������s���2��B��ɟ��3-F�������"��<����m�MC���m��<����"�����3-F�ɟ���B����2���s����`   `   �� �P����%���w�l�!�6�ʿv�v�%[�������@��ܽ���sN^�����ܽ��@�����%[�v�v�6�ʿl�!��w��%��P���`   `   �<�q�)�r���y
���!I��A���i����)�`�¾�?[����ث���@u�ث������?[�`�¾��)��i���A���!I�y
��r���q�)�`   `   �`o�$7W���-�����g�o�	�3M����:��WԾ��m�c�g��0]��g��c���m��WԾ��:�3M��o�	���g�-�����$7W�`   `   ڠ��Bi�S�)��4����s��u�Ҋ���^A�+�۾	�u��X	�襽섽襽�X	�	�u�+�۾�^A�Ҋ���u���s��4��S�)�Bi�`   `   O_o��:W��"�����h�-=
���,�<��z׾*�q�����/������/�����*�q��z׾,�<���-=
��h�����"��:W�`   `   -�<�S�)������r��"HJ�����Kؓ���-��>Ⱦ%�a�!7��y��� p�y���!7��%�a��>Ⱦ��-�Kؓ�����"HJ��r������S�)�`   `   w ��v���I��~x�t�"�a�ͿĽ|��X���[uH�-G�rn��	S�qn��-G�[uH����X�Ľ|�a�Ϳt�"�~x��I���v��`   `   y
��zI����s�]~3�{����ơ��dL�2��� ���c)�>s��P6_�$/�P6_�>s���c)�� ��2���dL��ơ�{���]~3���s�zI��`   `   �3L�5O@���!�����d��F,r��^�ִľkl��H�����\0�A���\0�����H�kl�ִľ�^�F,r��d�������!�5O@�`   `   �s ��A����ҿ���Tx���-������Mu4��_ѽ8_h�=h�Oʼ=h�8_h��_ѽMu4�����羞�-�Tx������ҿ�A��`   `   �`��(��������[��z'�.�������V�d�;��+�,���ü�ʔ���ü+�,�;��d��V�����.��z'���[�����(��`   `   &,F��>�j�)�1���۾����M�a�o�������+d�/��������~�����/���+d�����o��M�a�������۾1�j�)��>�`   `   O��v�SGҾ�^���֌�8�S����н�/��ۢ4�A��g���؍��g���A��ۢ4��/���н��8�S��֌��^��SGҾ�v�`   `   V���t��[&��(Q[���1��t	��wͽ�1���*a�I]/���q���j �q����I]/��*a��1���wͽ�t	���1�(Q[�[&��t��`   `   r�-�?�(�������Ӓ�P"�������_�)�f�y_���a���f��&i���f���a�y_�)�f��_�����P"��Ӓὰ�����?�(�`   `   �ν�ɽmY��P�����Kb���-��/ŉ�
3��!'��Ɨ��<̽yoѽ<̽Ɨ��!'��
3��/ŉ��-��Kb�����P��mY���ɽ`   `   �M|��y���q��Vk��>n�[)��z��������_佡Q
�*� ��=0�6�5��=0�*� ��Q
��_佇���z���[)���>n��Vk���q��y�`   `   z&�*c(�Z)0�M�C�z#k�䗽�&̽�w	��84�4�a����o��>G��o�����4�a��84��w	��&̽䗽z#k�M�C�Z)0�*c(�`   `   ���X��{����J�h����Tͽ����0R�R�>d���tپ��ke�����tپ>d��R��0R�����Tͽh�����J�{��X��`   `   '�鼑� ��](�\�u��]���Q�BW[�S5����۾��$�-�e6D��gL�e6D�$�-�����۾S5��BW[��Q��]��\�u��](��� �`   `   x���_���I�����xD �q�L��ʞ����m&�Z]�!݈��_��i����_��!݈�Z]�m&���뾘ʞ�q�L�xD ������I�_��`   `   4���A(��^{�A�ν/K,����ww߾w�)���u�1���dԿ�����������dԿ1�����u�w�)�ww߾���/K,�A�ν�^{��A(�`   `   p�'�FI�������q�`�1�����/�l��d��$J���_"�/JA��jM�/JA��_"�$J���d��/�l���1���q�`�������FI�`   `   MC���m��<����"�����3-F�ɟ���B����2���s����as�������s���2��B��ɟ��3-F�������"��<����m�`   `   sN^�����ܽ��@�����%[�v�v�6�ʿl�!��w��%��P����� �P����%���w�l�!�6�ʿv�v�%[�������@��ܽ���`   `   �@u�ث������?[�`�¾��)��i���A���!I�y
��r���q�)��<�q�)�r���y
���!I��A���i����)�`�¾�?[����ث��`   `   0]��g��c���m��WԾ��:�3M��o�	���g�-�����$7W��`o�$7W���-�����g�o�	�3M����:��WԾ��m�c�g��`   `   섽襽�X	�	�u�+�۾�^A�Ҋ���u���s��4��S�)�Bi�ڠ��Bi�S�)��4����s��u�Ҋ���^A�+�۾	�u��X	�襽`   `   ����/�����*�q��z׾,�<���-=
��h�����"��:W�O_o��:W��"�����h�-=
���,�<��z׾*�q�����/��`   `    p�y���!7��%�a��>Ⱦ��-�Kؓ�����"HJ��r������S�)�-�<�S�)������r��"HJ�����Kؓ���-��>Ⱦ%�a�!7��y���`   `   	S�qn��,G�[uH����X�Ľ|�a�Ϳt�"�~x��I���v��w ��v���I��~x�t�"�a�ͿĽ|��X���[uH�,G�qn��`   `   #/�P6_�=s���c)�� ��2���dL��ơ�{���]~3���s�zI��y
��zI����s�]~3�{����ơ��dL�2��� ���c)�=s��P6_�`   `   @���\0�����H�
kl�ִľ�^�F,r��d�������!�5O@��3L�5O@���!�����d��F,r��^�ִľ
kl��H�����\0�`   `   Nʼ<h�7_h��_ѽMu4�����羞�-�Tx������ҿ�A���s ��A����ҿ���Tx���-������Mu4��_ѽ7_h�<h�`   `   �ʔ���ü+�,�;��d��V�����.��z'���[�����(���`��(��������[��z'�.�������V�d�;��+�,���ü`   `   B��ù�/���4���Խ��'���|��s���������@���X���a���X��@��������s����|���'��Խ�4��/��ù�`   `   �
��b`˼޸
�� O�:�����.,�.[p�m쟾9�ɾ[R�@����	�@��[R�9�ɾl쟾.[p�.,���;���� O�޸
�b`˼`   `   �A����
v(��K�󺃽�>��I��Es �(�N���~�Ϫ��i|��Ш�i|��Ϫ����~�(�N�Es �I���>�������K�
v(����`   `   �����쀽�d�?�z����L��_,����὎$
�Ǘ$��.<��L�iwR��L��.<�Ǘ$��$
����_,���L��z���?��d��쀽`   `   �@罈�QԽ�����?������ x���E��\�Ƚ�G⽄o�����N		�����o���G�\�Ƚ�E�� x�������?������QԽ��`   `   �H���B�Up2�Z���t��ܽE8���ǭ�D۩�����h���\���7���\��h������D۩��ǭ�E8���ܽ�t�Z��Up2���B�`   `   (ĩ���5a��>�|�6�L�Av ��[��ɽ�t���#���\���䗽�'���䗽�\���#���t��ɽ�[��Av �6�L�>�|�5a����`   `   Y��ʫ����R˾T���q���0�J��Tǽf]�� Ð�죈��t��죈� Ð�f]���TǽJ���0��q�T��R˾���ʫ�`   `   ��f��i]���C�>� �1���2޴�w�~��1��w��%��9䗽�����������9䗽%���w���1�w�~�2޴�1���>� ���C��i]�`   `   K����"���-��{� W<�A������Jr���!�&��Ϩ�u)����u)��Ϩ�&����!�Jr�����A�� W<�{��-���"��`   `   e��V���������F����@�Dz��p�����P�A		�Rt��'ؗ�����'ؗ�Rt��A		���P�p���Dz����@��F����������V�`   `   ��x���h�L7A�Gq�]�˿�7����,��׾ő��&��vܽ�ߤ��0���ߤ��vܽ&�ő���׾��,��7��]�˿Gq�L7A���h�`   `   fL��f���{���`V���������a�`���|��g�E�(Z����������(Z��g�E��|��`����a��������`V��{��f��`   `   �.�����9��e��_W@�Ra����l\&�d¾�Rd�����.���֤��.������Rd�d¾l\&����Ra�_W@�e���9�����`   `   1U���h�.m)�X���Վs��
㦿��@��dݾ��~�,a�Q�Ƚ�A��Q�Ƚ,a���~��dݾ��@�
㦿�Վs�X���.m)��h�`   `   ������"�V�gL �|S���"�4���[�S�\E��V���� yͽ�Ϋ� yͽ���V��\E�[�S�4����"�|S��gL �"�V����`   `   ���6֟��h�Z5
�D{��f)������%[�A����z��>Z ��u˽�<���u˽>Z ��z��A����%[�����f)�D{��Z5
��h�6֟�`   `   ������5�V�#n �R�����"��Ӻ��yU�c����������p؞����������c���yU��Ӻ���"�R���#n �5�V����`   `   �O���h�F�)��K����t�V�����C�o�߾~�|�pW�����͏����pW�~�|�o�߾�C����V���t��K��F�)��h�`   `   ��-����`������M�A��h�p�����)�rľ�_�����F3���Ux�F3�������_�rľ��)�p����h�M�A�����`�����`   `   I���䖾�h{���W�gV������f�������8�;��ӽ�G��sK��G��ӽ8�;���������f����gV��W�h{��䖾�`   `   S�w���g���@������Ϳ����ې0�j�ھk���h���E��T~H����T~H��E��h��k���j�ھې0�������Ϳ�����@���g�`   `   A����wG�������X����C��}�P��k-G�3�<k��Wz��:�Wz�<k��3�k-G�P���}���C��X������wG����`   `   ����2���샚��z��=����N��Aim�����3sA�9༿��9�3sA�����Aim��N�����=��z�샚�2���`   `   ��a���X��@��������s����|���'��Խ�4��0��ù�B��ù�0���4���Խ��'���|��s���������@���X�`   `   ��	�@��[R�9�ɾm쟾.[p�.,���;���� O�޸
�c`˼�
��c`˼޸
�� O�;�����.,�.[p�m쟾9�ɾ[R�@��`   `   Ш�i|��Ϫ����~�(�N�Es �I���>�������K�
v(�����A����
v(��K������>��I��Es �(�N���~�Ϫ��i|��`   `   iwR��L��.<�Ǘ$��$
����_,���L��{���?��d��쀽�����쀽�d�?�{����L��_,����὎$
�Ǘ$��.<��L�`   `   O		�����o���G�]�Ƚ�E�� x�������?������QԽ�⽑@罈�QԽ�����?������ x���E��]�Ƚ�G⽄o�����`   `   �7���\��h������D۩��ǭ�F8���ܽ�t�Z��Up2���B��H���B�Up2�Z���t��ܽF8���ǭ�D۩�����h���\��`   `   �'���䗽�\���#���t��ɽ�[��Av �6�L�>�|�5a����(ĩ���5a��>�|�6�L�Av ��[��ɽ�t���#���\���䗽`   `   �t��죈� Ð�f]���TǽJ���0��q�T��R˾���ʫ�Y��ʫ����R˾T���q���0�J��Tǽf]�� Ð�죈�`   `   �������9䗽&���w���1�w�~�2޴�1���>� ���C��i]���f��i]���C�>� �1���2޴�w�~��1��w��%��9䗽����`   `   ��u)��Ϩ�&����!�Jr�����A�� W<�{��-���"��K����"���-��{� W<�A������Jr���!�&��Ϩ�u)��`   `   ����'ؗ�Rt��A		���P�p���Dz����@��F����������V�e��V���������F����@�Dz��p�����P�A		�Rt��'ؗ�`   `   �0���ߤ��vܽ&�ő���׾��,��7��]�˿Gq�L7A���h���x���h�L7A�Gq�]�˿�7����,��׾ő��&��vܽ�ߤ�`   `   �����(Z��g�E��|��`����a��������`V��{��f��fL��f���{���`V���������a�`���|��g�E�(Z�����`   `   �֤��.������Rd�d¾l\&����Ra�_W@�e���9������.�����9��e��_W@�Ra����l\&�d¾�Rd�����.��`   `   �A��P�Ƚ,a���~��dݾ��@�
㦿�Վs�Y���.m)��h�1U���h�.m)�X���Վs��
㦿��@��dݾ��~�,a�P�Ƚ`   `   �Ϋ� yͽ���V��\E�[�S�4����"�}S��gL �"�V����������"�V�gL �|S���"�4���[�S�\E��V���� yͽ`   `   �<���u˽>Z ��z��A����%[�����f)�D{��Z5
��h�6֟����6֟��h�Z5
�D{��f)������%[�@����z��>Z ��u˽`   `   o؞����������c���yU��Ӻ���"�R���#n �5�V����������5�V�#n �R�����"��Ӻ��yU�c����������`   `   �͏����pW�~�|�o�߾�C����V���t��K��F�)��h��O���h�F�)��K����t�V�����C�o�߾~�|�pW����`   `   �Ux�F3�������_�rľ��)�p����h�M�A�����`�������-����`������M�A��h�p�����)�rľ�_�����F3��`   `   �sK��G��ӽ8�;���������f����gV��W�h{��䖾�I���䖾�h{���W�gV������f�������8�;��ӽ�G�`   `   ���S~H��E��h��k���j�ھې0�������Ϳ�����@���g�S�w���g���@������Ϳ����ې0�j�ھk���h���E��S~H�`   `   �:�Vz�<k��3�k-G�P���}���C��X������vG����A����vG�������X����C��}�P��k-G�3�<k��Vz�`   `   ���9�3sA�����Aim��N�����=��z�샚�2�������2���샚��z��=����N��Aim�����3sA�9�`   `   #ߢ���ɼ�"�(��x��>�1�I���fͿ����j�(���K��je�Y�n��je���K�j�(����fͿ�I���>�1�x��(���"���ɼ`   `   �:ü-Lݼ���!c�����/�~;��	���s����ؾ_| �y��F��y��_| ���ؾ�s���	��~;��/�����!c���-Lݼ`   `   ���"���8�9d��l��q�ɽ��:v5�F�h��x��}���ڰ��tu��ڰ��}����x��F�h�:v5���r�ɽ�l��9d���8��"�`   `   �|������Q��sŏ�������]�ݽG��S�&�S_E�<�`��@s�n�y��@s�<�`�S_E�S�&�G��]�ݽ������sŏ�Q������`   `   D���y���ӽ��ɽR�Ƚ�ӽ�l�nS�Z��B�%���0���4���0�B�%�Z��nS��l��ӽR�Ƚ��ɽ�ӽy�Ὢ��`   `   6NP�.�J�W�;���&����h� �������L𽁫���X���%6����X������L𽯱轌��h� ������&�W�;�.�J�`   `   ���0j��!��d��� �]��x5�+�EV�`f������Y������� �����Y�����`f��EV�+��x5� �]�d���!��0j��`   `   �T�m��8���Bվu����p��H�L�)�#��j�Y���)v���	��*3���	��)v��Y����j�)�#�H�L��p��u����Bվ�8��m�`   `   +�p�V�f�a�L��(�G��O�¾i}����S�2�%� ����� ��ʦ� ����� �2�%���S�i}��O�¾G���(�a�L�V�f�`   `   �Ŀ6ݻ�ﱣ�����,.F�� ��zƾ�芾�J�J$�C!�k~��0��k~��C!�J$��J��芾�zƾ� �,.F�����ﱣ�6ݻ�`   `   8!�f��P�r�ʿ����b�K�o������Hx�$�4�ޘ�$��d?��$��ޘ�$�4�Hx�����o��b�K�����r�ʿP�f��`   `   F^��/y�C�M�����ֿ2���z�7�$�龈����"O�^��&�t����&�^��"O�����$��z�7�2����ֿ���C�M�/y�`   `   �f������������d�U��[���	�n�������i5k�?�%��#�5����#�?�%�i5k�������	�n�[���U����d���������`   `   �aA�.�x �h����L�۽���ɔ�y�0�X�Ӿ_-���,/��
�=1��
��,/�_-��X�Ӿy�0��ɔ�۽����L�h��x �.�`   `   6܏��a���A<�����f������ޯ��K����gu��P6�8B�=�8B�P6�gu������K��ޯ���f��������A<��a��`   `   �~��\(���n����h����+�osÿI�^�����|��p�8��S2��p�8��|�����I�^�osÿ��+�h������n�\(��`   `   D,��ٴ���a���T�����3� �ʿ�f����ة��lb5�����ҽ���lb5�ة������f� �ʿ��3�T�����a��ٴ��`   `   ~��N*��D�n��������I�,��MĿ�_����`@����+����4߿������+�`@������_��MĿI�,��������D�n�N*��`   `   ׏��a��}Z<�4f��{��؎��C��B�L�꾑���G���ɽ|v����ɽG������B�L��C��؎�{��4f��}Z<��a��`   `   'EA��.��� ����]N����8��"�0��̾�ij�f���
���ۍ��
��f���ij��̾"�0��8����]N������ ��.�`   `   �����6��J���d�e����x�¿n�p�}���f��D�0jὴ��P�c����0j�D��f��}��n�p�x�¿���d�e�J����6��`   `   �̄�pGx��OM��B��ؿ}ɏ���7�7��x�����qֲ�,<Y���-�,<Y�qֲ����x��7����7�}ɏ��ؿ�B��OM�pGx�`   `   O��I������ʿ�$��نL�����i����N�f�As��r�!�`���r�!�As��f���N��i�����نL��$���ʿ���I��`   `   �¿��������c���OF�0Q�&���ux�M�����M����q������M����M�ux�&���0Q��OF��c���������`   `   Y�n��je���K�j�(����fͿ�I���>�1�x��(���"���ɼ$ߢ���ɼ�"�(��x��>�1�I���fͿ����j�(���K��je�`   `   F��y��_| ���ؾ�s���	��~;��/�����!c���-Lݼ�:ü-Lݼ���!c�����/�~;��	���s����ؾ_| �y��`   `   uu��ڰ��}����x��F�h�:v5���r�ɽ�l��9d���8��"����"���8�9d��l��r�ɽ��:v5�F�h��x��}���ڰ��`   `   n�y��@s�<�`�S_E�S�&�G��]�ݽ������sŏ�Q�������|������Q��sŏ�������]�ݽG��S�&�S_E�<�`��@s�`   `   ��4���0�C�%�Z��nS��l��ӽR�Ƚ��ɽ�ӽy�Ὢ��D���y���ӽ��ɽR�Ƚ�ӽ�l�nS�Z��C�%���0�`   `   %6����X������L𽯱轌��h� ������&�W�;�.�J�6NP�.�J�W�;���&����h� �������L𽁫���X���`   `   �� �����Y�����af��EV�+��x5� �]�d���!��0j�����0j��!��d��� �]��x5�+�EV�`f������Y�����`   `   *3���	��)v��Y����j�)�#�I�L��p��u����Bվ�8��m��T�m��8���Bվu����p��H�L�)�#��j�Y���)v���	��`   `   ˦� ����� �2�%���S�i}��O�¾G���(�a�L�V�f�+�p�V�f�a�L��(�G��O�¾i}����S�2�%� ����� ��`   `   0��l~��D!�J$��J��芾�zƾ� �-.F�����ﱣ�6ݻ��Ŀ6ݻ�ﱣ�����,.F�� ��zƾ�芾�J�J$�D!�l~��`   `   d?��$��ޘ�$�4�Hx�����o��b�K�����r�ʿP�f��8!�f��P�r�ʿ����b�K�o������Hx�$�4�ޘ�$��`   `   t����&�^��"O�����$��{�7�2����ֿ���C�M�/y�F^��/y�C�M�����ֿ2���z�7�$�龈����"O�^��&�`   `   5����#�?�%�i5k�������	�n�[���U����d����������f������������d�U��[���	�n�������i5k�?�%��#�`   `   =1��
��,/�_-��X�Ӿy�0��ɔ�۽����L�h���x �.��aA�.�x �h����L�۽���ɔ�y�0�X�Ӿ_-���,/��
�`   `   =�8B�P6�gu������K��ޯ���f��������A<��a��6܏��a���A<�����f������ޯ��K����gu��P6�8B�`   `   S2��p�8��|�����I�^�osÿ��+�h������n�\(���~��\(���n����h����+�osÿI�^�����|��p�8��`   `   �ҽ���lb5�ة������f� �ʿ��3�T�����a��ٴ��D,��ٴ���a���T�����3� �ʿ�f����ة��lb5����`   `   4߿������+�`@������_��MĿI�,��������D�n�N*��~��N*��D�n��������I�,��MĿ�_����`@����+����`   `   |v����ɽG������B�L��C��؎�{��4f��}Z<��a��׏��a��}Z<�4f��{��؎��C��B�L�꾑���G���ɽ`   `   �ۍ��
��f���ij��̾"�0��8����]N������ ��.�'EA��.��� ����]N����8��"�0��̾�ij�f���
��`   `   P�c����0j�D��f��}��n�p�x�¿���d�e�J����6�������6��J���d�e����x�¿n�p�}���f��D�0jέ��`   `   ��-�+<Y�qֲ����x��7����7�}ɏ��ؿ�B��OM�pGx��̄�pGx��OM��B��ؿ}ɏ���7�7��x�����qֲ�+<Y�`   `   _���q�!�As��f���N��i�����نL��$���ʿ���I��O��I������ʿ�$��نL�����i����N�f�As��q�!�`   `   q������M����M�ux�&���/Q��OF��c����������¿��������c���OF�/Q�&���ux�M�����M����`   `   a��i\ּg*�c:��\�罬5�r.�����8��tq'�+�I�~Pb��\k�~Pb�+�I�tq'�8�����r.���5�\��c:��g*�i\ּ`   `   �:ϼA켤_#�x'u��͹���	�e�E�27��K����߾H���������H����߾K��27��e�E���	��͹�x'u��_#�A�`   `    � ��*��;G�h�|�󩨽��k��5K�������������kž�b˾�kž������������5K�k���󩨽h�|��;G��*�`   `   �c������4͑�<�������/5ڽi��g&�`@J�x0n�����&:������&:������x0n�`@J�g&�i��/5ڽ����<���4͑�����`   `   ��q����罰0���b��;�#O���0�j.I�ٗ^�Em��~r�Em�ٗ^�j.I���0�#O�;�b���影0����q��`   `   T�L��XH�ȑ<�JW-��{������N���a+���;�
K���U���Y���U�
K���;��a+�N��������{�JW-�ȑ<��XH�`   `   &�������JF��?-���mi�.7K��8�{�0�|l3��&<���F���N���Q���N���F��&<�|l3�{�0��8�.7K��mi�?-��JF������`   `   ������p����Ӿ�:�������l���P�E��}D��GI��iN���P��iN��GI��}D�E���P��l������:����Ӿ�p�����`   `   =�g���^�_$F��$�h���xɾ+����~�8�^��HQ���N�}�O���P�}�O���N��HQ�8�^��~�+����xɾh���$�_$F���^�`   `   z��� ���n��m�O�B��6��jѾx�����A�`��1T�krP���O�krP��1T�A�`����x���jѾ�6�O�B�m��n��� ��`   `   �����L��h�¿�C��H�I�r���rž���x�r���X���N��L���N���X�x�r�����ržr��H�I��C��h�¿�L����`   `   3z�U-j�h`B���ܖο�(����7��/��쭫��ۂ��o\�NNJ��XE�NNJ��o\��ۂ�쭫��/����7��(��ܖο��h`B�U-j�`   `   US��m߿�8S����W�ԏ�W2���ak���&qžp����^�Z�C��<�Z�C��^�p���&qž���ak�W2��ԏ���W�8S��m߿�`   `   ��.����o��V ��F�A�
���/1�1�޾YÕ�v�^�/,;���0�/,;�v�^�YÕ�1�޾/1����
��F�A�V ���o����`   `   Eځ�A�i�$9*���O>u����=@��b�I����u���sz\�7�0��$�7�0�sz\�u������b�I�=@�����O>u���$9*�A�i�`   `   ~����7��x�W��� �R2��Th#�FL����Z�V/�����9V��P$�����P$��9V����V/���Z�FL��Th#�R2���� �x�W��7��`   `   &O���o��$�i���
��R����*���¿�3`���R ��)K�8�����8��)K�R �����3`���¿��*��R����
�$�i��o��`   `   Ӹ��y9����W����k����#�b\����X�ek��ߔ���:�����������:�ߔ�ek����X�b\����#��k������W�y9��`   `   �Ձ��i�M*��R����u���^��4$F��2�^)����%�%�佄ƽ%����%�^)���2�4$F�^������u��R��M*��i�`   `   y�.����f����O���B��p￾O���+���Ⱦ��j����ս�G���ս������j���Ⱦ�+��O���p��B��O��f������`   `   ���P����R��pGX���MO���g�6j�T���w(C���罛��2�|�������w(C�T���6j��g�MO����pGX��R��P���`   `   �Ry���i��+B������ο�N��4�1��Lܾ󐄾����7���Jf��<��Jf��7�����󐄾�Lܾ4�1��N����ο����+B���i�`   `   t�\��������¿7쎿�$F� �W���"�K���{���t*�j�t*�{�����"�K�W��� ��$F�7쎿��¿����\��`   `   �O��n���.���=��5�A���
��鼾��u�l$�Xa��LnR������Jɼ����LnR�Xa��l$���u��鼾��
�5�A�=��.���n���`   `   �\k�~Pb�+�I�tq'�8�����r.���5�\��c:��g*�j\ּa��j\ּg*�c:��\�罬5�r.�����8��tq'�+�I�~Pb�`   `   �����H����߾K��27��e�E���	��͹�x'u��_#�A켛:ϼA켤_#�x'u��͹���	�e�E�27��K����߾H����`   `   �b˾�kž������������5K�k���󩨽h�|��;G��*� � ��*��;G�h�|�󩨽��k��5K�������������kž`   `   ����&:������x0n�`@J�g&�i��/5ڽ����<���4͑������c������4͑�<�������/5ڽi��g&�`@J�x0n�����&:��`   `   �~r�Em�ٗ^�j.I���0�#O�;�c���影0����q����q����罱0���c��;�#O���0�j.I�ٗ^�Em�`   `   ��Y���U�
K���;��a+�N��������{�JW-�ȑ<��XH�T�L��XH�ȑ<�JW-��{������N���a+���;�
K���U�`   `   ��Q���N���F��&<�|l3�{�0��8�.7K��mi�?-��JF������&�������JF��?-���mi�.7K��8�{�0�|l3��&<���F���N�`   `   ��P��iN��GI��}D�E���P��l������:����Ӿ�p�����������p����Ӿ�:�������l���P�E��}D��GI��iN�`   `   ��P�}�O���N��HQ�8�^��~�+����xɾh���$�_$F���^�=�g���^�_$F��$�h���xɾ+����~�8�^��HQ���N�}�O�`   `   ��O�krP��1T�A�`����x���jѾ�6�O�B�m��n��� ��z��� ���n��m�O�B��6��jѾx�����A�`��1T�krP�`   `   �L���N���X�x�r�����ržr��H�I��C��h�¿�L���������L��h�¿�C��H�I�r���rž���x�r���X���N�`   `   �XE�NNJ��o\��ۂ�쭫��/����7��(��ܖο��h`B�U-j�3z�U-j�h`B���ܖο�(����7��/��쭫��ۂ��o\�NNJ�`   `   �<�Z�C��^�p���&qž���ak�W2��ԏ���W�8S��m߿�US��m߿�8S����W�ԏ�W2���ak���&qžp����^�Z�C�`   `   ��0�/,;�v�^�YÕ�1�޾/1����
��F�A�V ���o������.����o��V ��F�A�
���/1�1�޾YÕ�v�^�/,;�`   `   �$�7�0�sz\�u������b�I�=@�����O>u���$9*�A�i�Eځ�A�i�$9*���O>u����=@��b�I����u���sz\�7�0�`   `   ����P$��9V����V/���Z�FL��Th#�R2���� �x�W��7��~����7��x�W��� �R2��Th#�FL����Z�V/�����9V��P$�`   `   ���8��)K�R �����3`���¿��*��R����
�$�i��o��&O���o��$�i���
��R����*���¿�3`���R ��)K�8��`   `   �������:�ߔ�ek����X�b\����#��k������W�y9��Ӹ��y9����W����k����#�b\����X�ek��ߔ���:����`   `   �ƽ%����%�^)���2�4$F�^������u��R��M*��i��Ձ��i�M*��R����u���^��4$F��2�^)����%�%��`   `   G���ս������j���Ⱦ�+��O���p��B��O��f������y�.����f����O���B��p￾O���+���Ⱦ��j����ս�`   `   2�|�������w(C�T���6j��g�MO����pGX��R��P������P����R��pGX���MO���g�6j�T���w(C���罛��`   `   �<��Jf��7�����󐄾�Lܾ4�1��N����ο����+B���i��Ry���i��+B������ο�N��4�1��Lܾ󐄾����7���Jf�`   `   j�s*�z�����"�K�W��� ��$F�7쎿��¿����\��t�\��������¿7쎿�$F� �W���"�K���z���t*�`   `   �Jɼ����KnR�Xa��l$���u��鼾��
�5�A�=��.���n����O��n���.���=��5�A���
��鼾��u�l$�Xa��KnR�����`   `   ݕ��8H��G4�j\����T5�6������,9�� ���s=��qS��x[��qS��s=� ��,9������6��T5���j\���G4�8H�`   `   KA�_� �3����'}ɽ���P��h��XG����(��!����!�(����XG���h���P���'}ɽ���3�_� �`   `   B(��C4��MZ����N½Dq���1�Kg��Ԑ��ӭ�s�ƾ�׾|�ݾ�׾s�ƾ�ӭ��Ԑ�Kg���1�Dq��N½���MZ��C4�`   `   ����e��F���&ű���ֽ���$�'�cP�Ǐ|��֓�"���u��oѶ��u��"���֓�Ǐ|�cP�$�'������ֽ&ű�F���e��`   `   l��轰��}���:o����5�.��WN�c�q�Ds���f��y��K��y���f��Ds��c�q��WN�5�.����:o�}��������`   `   �A���>�Is8�g(2�t�/��I5�Q�C���Z�:pw�\���%ܗ��ؠ�
���ؠ�%ܗ�\���:pw���Z�Q�C��I5�t�/�g(2�Is8���>�`   `   /e���Κ�	L����+,t�9g�Lf���q�IJ��cƏ�Bw��涣�Ѯ��涣�Bw��cƏ�IJ����q�Lf�9g�+,t���	L���Κ�`   `   �� ��y��^���"ɾ�����;��
���'툾�����z���7��:����:��:����7���z������'툾
����;�������"ɾ^�侗y��`   `   � O�P�G�Wm3�#r�x:��G�̾ح�����bj�����Z���>����̫�>���Z������bj������ح�G�̾x:��#r�Wm3�P�G�`   `   �p��)t��^Ӌ��Jf�J�4��W�s۾����Ħ�����Ф��a�������a���Ф�����Ħ����s۾�W�J�4��Jf�^Ӌ�)t��`   `   �i�����R�׿�D��즁��w=�ku�.�׾ɽ������=������0X�������=�����ɽ��.�׾ku��w=�즁��D��R�׿����`   `   �O��C��$��z���۶�9m~�pz0��W��WƾM����G���蛾FZ���蛾�G��M���Wƾ�W��pz0�9m~��۶��z���$��C�`   `   �K��Z��r-w��5�)���팦�G[������׾6���h��O���ŏ�O����h��6����׾���G[�팦�)����5�r-w�Z��`   `   ��[(���R��6{��$���ѿ�a���~*���ڑ������Ʌ����Ʌ����ڑ���辏~*��a����ѿ�$�6{��R��[(��`   `   ya>�@|+�?����&����L�#����똿qx=����&׭�{J��Q�q�m�h�Q�q�|J��&׭����qx=��똿#�����L��&��?���@|+�`   `   Ƃq�6Y���G+��<Qk��]�k_��I�I�����i�=T~���V��K���V�=T~�i񩾐���I�I�k_���]�<Qk�G+����6Y�`   `   :���O0k�'|+�Z���U-w����E����L�g<��9򡾲g�8Y;�y�.�8Y;��g�9�g<����L�E�����U-w�Z���'|+�O0k�`   `   Łq�"8Y�ʻ�CE��bsk��:�e(���E��}�I����L�����j�����L�I����}��E�e(���:�bsk�CE��ʻ�"8Y�`   `   �[>��{+�)���iK����L�3����J��No3�c׾X���G0�.i���.i��G0�X��c׾No3��J��3�����L�iK��)����{+�`   `   )�����[`��!k{�H�$��п���F �
���&�c���0�ԽK��0�Խ��&�c�
���F �����пH�$�!k{�[`�����`   `   �%���@��,w���5�����&���O�Q9���њ���;��뽥���% �������뽡�;��њ�Q9��O�&���������5�,w��@��`   `   ��O�"�C�{�$�A���]��0-v�S= �޼ɾ�hw�^{�s=��U2v�Q�U2v�s=��^{��hw�޼ɾS= �0-v��]��A��{�$�"�C�`   `   8��f�����ؿC��5��wn3�Is�Қ�}s@�@r�����<4��^��<4����@r�}s@��Қ�Is�wn3�5��C����ؿf���`   `   �X��%@��}!��bh���1�j� ��㱾��j�3���ڴ�[QW�Θ�J�ܼΘ�[QW��ڴ�3����j��㱾j� ���1�bh�}!��%@��`   `   �x[��qS��s=� ��,9������6��T5���j\���G4�8H�ݕ��8H��G4�j\����T5�6������,9�� ���s=��qS�`   `   ���!�(����XG���h���P���'}ɽ���3�`� �KA�`� �3����'}ɽ���P��h��XG����(��!�`   `   |�ݾ�׾s�ƾ�ӭ��Ԑ�Kg���1�Dq��N½���MZ��C4�B(��C4��MZ����N½Dq���1�Kg��Ԑ��ӭ�s�ƾ�׾`   `   oѶ��u��"���֓�Ǐ|�cP�$�'������ֽ&ű�F���e������e��F���&ű���ֽ���$�'�cP�Ǐ|��֓�"���u��`   `   L��y���f��Ds��c�q��WN�6�.����:o�}��������l��轰��}���:o����6�.��WN�c�q�Ds���f��y��`   `   
���ؠ�%ܗ�\���:pw���Z�Q�C��I5�t�/�g(2�Is8���>��A���>�Is8�g(2�t�/��I5�Q�C���Z�:pw�\���%ܗ��ؠ�`   `   Ѯ��涣�Bw��cƏ�IJ����q�Lf�9g�+,t���	L���Κ�/e���Κ�	L����+,t�9g�Lf���q�IJ��cƏ�Bw��涣�`   `   �:��:����7���z������'툾
����;�������"ɾ^�侗y���� ��y��^���"ɾ�����;��
���'툾�����z���7��:���`   `   �̫�>���Z������bj������ح�G�̾x:��#r�Wm3�P�G�� O�P�G�Wm3�#r�x:��G�̾ح�����bj�����Z���>���`   `   �����a���Ф�����Ħ����s۾�W�J�4��Jf�^Ӌ�)t���p��)t��^Ӌ��Jf�J�4��W�s۾����Ħ�����Ф��a��`   `   0X�������=�����ɽ��.�׾ku��w=�즁��D��R�׿�����i�����R�׿�D��즁��w=�ku�.�׾ɽ������=������`   `   FZ���蛾�G��M���Wƾ�W��pz0�9m~��۶��z���$��C��O��C��$��z���۶�9m~�pz0��W��WƾM����G���蛾`   `   ŏ�O����h��6����׾���G[��)����5�r-w�Z���K��Z��r-w��5�)���팦�G[������׾6���h��O���`   `   ���Ʌ����ڑ���辏~*��a����ѿ�$�6{��R��[(����[(���R��6{��$���ѿ�a���~*���ڑ������Ʌ�`   `   m�h�Q�q�|J��&׭����rx=��똿#�����L��&��?���@|+�ya>�@|+�?����&����L�#����똿qx=����&׭�{J��Q�q�`   `   �K���V�=T~�i񩾐���I�I�k_���]�<Qk�G+����6Y�Ƃq�6Y���G+��<Qk��]�k_��I�I�����i�=T~���V�`   `   y�.�8Y;��g�9�g<����L�E�����U-w�Z���'|+�O0k�:���O0k�'|+�Z���U-w����E����L�g<��9򡾲g�8Y;�`   `   �j�����L�I����}��E�e(���:�bsk�CE��ʻ�"8Y�Łq�"8Y�ʻ�CE��bsk��:�e(���E��}�I����L����`   `   ��.i��G0�X��c׾No3��J��3�����L�iK��)����{+��[>��{+�)���iK����L�3����J��No3�c׾X���G0�.i�`   `   K��0�Խ��&�c�
���F �����пH�$�!k{�[`�����)�����[`��!k{�H�$��п���F �
���&�c���0�Խ`   `   % �������뽡�;��њ�Q9��O�&���������5�,w��@���%���@��,w���5�����&���O�Q9���њ���;��뽤���`   `   Q�T2v�s=��^{��hw�޼ɾS= �0-v��]��A��{�$�"�C���O�"�C�{�$�A���]��0-v�S= �޼ɾ�hw�^{�s=��T2v�`   `   �^��<4����@r�}s@��Қ�Is�wn3�5��C����ؿf���8��f�����ؿC��5��wn3�Is�Қ�}s@�@r�����<4�`   `   J�ܼ͘�[QW��ڴ�3����j��㱾j� ���1�bh�}!��$@���X��$@��}!��bh���1�j� ��㱾��j�3���ڴ�[QW�͘�`   `   �8㼂x��-G�윽O��B�6�P���B��Ɵ쾾����-�΂@�>G�΂@���-����Ɵ쾙B��P��B�6�O��윽�-G��x�`   `   ���S`�B\M��T��ݴίz"��Aa�H֕�{���2��w��:��%�:��w��2��{���H֕��Aa��z"�ݴὅT��B\M�S`�`   `   �6��#G�fby�GT���I轏��`�S�UA��̨�vUȾ(�����q�����(�vUȾ̨�UA��`�S�����I�GT��fby��#G�`   `   �r���9���V����ν}P�
)���W�����)����达��վ�徶t��徉�վ�达)���������W�
)�}P���ν�V���9��`   `   �}���佮����)���p?�i�i�F����騾��¾)�ؾ5.�8H�5.�)�ؾ��¾�騾F���i�i��p?�)����������`   `   �L2�`|2��/4�g[:�I�H��ta�u������ٜ;�e�8��+��8�e�ٜ;������u�ta�I�H�g[:��/4�`|2�`   `   ���#B��������/���l@��:��n꨾f���ھ�ﾳ������������ھf��n꨾:��l@��/���������#B��`   `   o�ݾ��ؾ��˾���*.��A)��2����Z��b�;���T���:���:�T������b�;�Z��2���A)��*.�������˾��ؾ`   `   ��-�l(��K���g���Ӿ�XȾ�"˾�ؾL��s����,�p���,�s���L���ؾ�"˾�XȾ�Ӿg�����K�l(�`   `   �񆿯ၿ��h��QE��"����!���޾K�ᾧ9]����������]���9�K����޾�!쾊��"��QE���h��ၿ`   `   ivϿ�Dƿ2������t_�B�-���4��] 龠M�}���ȶ����ȶ��}����M�] �4����B�-��t_����2���Dƿ`   `   37�������ʿ��!U_�,�'��>�,����32��5��|��5�32���,�ﾀ>�,�'�!U_����ʿ�����`   `   /�i�ci[���7�[D�/�ɿj���KEG���W���޾��ؾ$8پCھ$8پ��ؾ�޾W����KEG�j���/�ɿ[D���7�ci[�`   `   @��H�����}�Qm:��� �Å��ĸg�Ų"��9��`Ծ��žt�������t�����ž`Ծ�9��Ų"�ĸg�Å���� �Qm:���}�H���`   `   ���ػ���ǥ���i������ɿ`D����-��o��\Ⱦ�����먾�֦��먾����\Ⱦ�o����-�`D����ɿ�����i��ǥ�ػ��`   `   ����J��-�������0�|�޿r���T:4�����ZX���������"2���������ZX������T:4�r���|�޿�0������-���J�`   `   �`��^�����������7�͸����4X3�M��p��XC���Hr���i��Hr�XC��p��M��4X3����͸忾�7����������^�`   `   ]���J��/��Ǭ����/���ܿ]ވ�7n*��d۾�u���g�2�F�%=�2�F��g��u���d۾7n*�]ވ���ܿ��/�Ǭ���/���J�`   `   ������Kƥ���i�T�7Fƿ��w��O��þ����D@����������D@�����þ�O���w�7FƿT���i�Kƥ����`   `   ���ߚ���}��:�{%��Z#����T�H��)����[�@9�����U�㽪���@9���[��)��H���T�Z#��{%���:��}�ߚ��`   `   ��i�k�[��7����1Eƿ����t�-�k�ܾI���3����㹽�T���㹽���3�I��k�ܾt�-�����1Eƿ����7�k�[�`   `   �������M ���ɿޓ��kM�A���ڰ�>T`��P��2��|����q�|���2���P�>T`��ڰ�A���kM�ޓ���ɿ�M ����`   `   X3ӿ�ɿyR��P~��)�W��M�r6Ӿ�H��S_2��� +���,G�}�+��,G� +����S_2��H��r6Ӿ�M�)�W�P~��yR���ɿ`   `   \d���ӈ�
hs�:�I��!�e��|����\�7���Q�� c��W�Ӗ ��W� c��Q��7����\��|��e��!�:�I�
hs��ӈ�`   `   >G�΂@���-����Ɵ쾚B��P��B�6�O��윽�-G��x��8㼂x��-G�윽O��B�6�P���B��Ɵ쾾����-�΂@�`   `   %�:��w��2��{���H֕��Aa��z"�޴ὅT��C\M�S`����S`�B\M��T��޴ίz"��Aa�H֕�{���2��w��:��`   `   �q�����(�vUȾ̨�UA��`�S�����I�GT��fby��#G��6��#G�fby�GT���I轏��`�S�UA��̨�vUȾ(����`   `   �t��徉�վ�达)���������W�
)�}P���ν�V���9���r���9���V����ν}P�
)���W�����)����达��վ��`   `   8H�5.�)�ؾ��¾�騾F���i�i��p?�)���������佟}���佮����)���p?�i�i�F����騾��¾)�ؾ5.�`   `   �+��8�e�ٜ;������u�ta�I�H�g[:��/4�`|2��L2�`|2��/4�g[:�I�H��ta�u������ٜ;�e�8�`   `   ���������ھf��n꨾:��l@��/���������#B�����#B��������/���l@��:��n꨾f���ھ�ﾳ���`   `   ��:�U������b�;�Z��2���A)��*.�������˾��ؾo�ݾ��ؾ��˾���*.��A)��2����Z��b�;���U���:�`   `   p���,�s���L���ؾ�"˾�XȾ�Ӿg�����K�l(���-�l(��K���g���Ӿ�XȾ�"˾�ؾL��s����,�`   `   ������]���9�K����޾�!쾊��"��QE���h��ၿ�񆿯ၿ��h��QE��"����!���޾K�ᾧ9]����`   `   ��ȶ��}����M�] �4����B�-��t_����2���DƿivϿ�Dƿ2������t_�B�-���4��] 龡M�}���ȶ��`   `   �|��5�32���,�ﾀ>�,�'�!U_����ʿ�����37�������ʿ��!U_�,�'��>�,����32��5�`   `   Cھ$8پ��ؾ�޾W����KEG�j���/�ɿ[D���7�ci[�/�i�ci[���7�[D�/�ɿj���KEG���W���޾��ؾ$8پ`   `   ����t�����ž`Ծ�9��Ų"�ĸg�Å���� �Qm:���}�H���@��H�����}�Qm:��� �Å��ĸg�Ų"��9��`Ծ��žt���`   `   �֦��먾����\Ⱦ�o����-�`D����ɿ�����i��ǥ�ػ�����ػ���ǥ���i������ɿ`D����-��o��\Ⱦ�����먾`   `   "2���������ZX������T:4�r���|�޿�0������-���J�����J��-�������0�|�޿r���T:4�����ZX���������`   `   ��i��Hr�XC��p��M��4X3����͸忾�7����������^��`��^�����������7�͸����4X3�M��p��XC���Hr�`   `   %=�2�F��g��u���d۾7n*�]ވ���ܿ��/�Ǭ���/���J�]���J��/��Ǭ����/���ܿ]ވ�7n*��d۾�u���g�2�F�`   `   ������D@�����þ�O���w�7FƿT���i�Kƥ����������Kƥ���i�T�7Fƿ��w��O��þ����D@����`   `   U�㽪���@9���[��)��H���T�Z#��{%���:��}�ߚ�����ߚ���}��:�z%��Z#����T�H��)����[�@9�����`   `   �T���㹽���3�I��k�ܾt�-�����1Eƿ����7�k�[���i�k�[��7����1Eƿ����t�-�k�ܾI���3����㹽`   `   ��q�|���2���P�>T`��ڰ�A���kM�ޓ���ɿ�M �����������M ���ɿޓ��kM�A���ڰ�>T`��P��2��|��`   `   }�+��,G��*����S_2��H��r6Ӿ�M�)�W�P~��yR���ɿX3ӿ�ɿyR��P~��)�W��M�r6Ӿ�H��S_2����*���,G�`   `   Ӗ ��W�c��Q��7����\��|��e��!�:�I�
hs��ӈ�\d���ӈ�
hs�:�I��!�e��|����\�7���Q��c��W�`   `   =G��<%���h��O���Q���>�M;��*������"��2���7��2��"���*���M;����>��Q��O����h��<%�`   `   �����5��Hx��`��	"���:��d~�g*��8�Ͼ���������������������8�Ͼg*���d~���:�	"��`���Hx���5�`   `   +�R��h�S����νG'�[�E��*���ݧ��lξ�B�
	��T�����T�
	��B�lξ�ݧ��*��[�E�G'��νS����h�`   `   �!��Mǡ��h½%����,&�v�[�����&�����ھ0^�������=�������0^����ھ&�������v�[��,&�%����h½Mǡ�`   `   �	߽-��@G����n�E��<{����X�žӃ�
�����m%�$)��m%������
�Ӄ�X�ž����<{�n�E����@G�-��`   `   �&�K�)�+&5��0K�>�n����Uj���AھQ��G�dh(�ů3�_�7�ů3�dh(�G�Q���AھUj�����>�n��0K�+&5�K�)�`   `   ڂx�;qy�r�}��4��!��Wۧ�oǾ���8�q�"���4�/P@��iD�/P@���4�q�"��8���oǾWۧ�!���4��r�}�;qy�`   `   lj������q`���ͱ��y��[-þ��ܾ2L �*����*��<��H�M��H��<���*�*��2L ���ܾ[-þ�y���ͱ�q`������`   `   ������ ]��1�E�S��cD���>��Q�.�Q@�uL��P�uL�Q@�Q�.�>����cD�S��E徙1� ]����`   `   *�P�!�J�>:�U%����k��&�.����-<.�<(>�`I��L�`I�<(>�-<.����.�&�k�����U%�>:�!�J�`   `   R��K�������b�o�=�Í"���mX�z���&)��6��Q@�C�C��Q@��6��&)�z��mX���Í"�o�=���b����K��`   `   $߿�6տ�X��o&��T�t�c�C�39%�e.��h�X ��v*�k\2� L5�k\2��v*�X ��h�e.�39%�c�C�T�t�o&���X���6տ`   `   ;������B ��r̿o]��n4j���7�ϻ��Y�{�����:t ���"�:t ����{���Y�ϻ���7�n4j�o]���r̿�B ����`   `   ��S�J�G��(�w���'C���[J�܏ �a����	�3�^��3�	����a�܏ ��[J�'C����w��(�J�G�`   `   R���^|�d�P�<���_�=^��Z��"����oK�{���ѥ��{�oK󾟥��"�Z�=^���_�<��d�P��^|�`   `   P����S���bp�_32��N��̴���Qc�G!�I���^�־��ɾoƾ�žoƾ��ɾ^�־I���G!��Qc�̴���N��_32��bp��S��`   `   �٧�Ԛ���^|���9�LC �8��&�b�dq�C&�򺾕㧾�Ƞ�� ���Ƞ��㧾�C&�dq�&�b�8��LC ���9��^|�Ԛ��`   `   χ���P���<p��1�f��,����W����!.;-���X���$��z��$�X��-���!.;�����W�,��f���1��<p��P��`   `   m����]|�4�P������ܿ�L���IC�Tc�~����?��v,[���E��{?���E�v,[��?��~���Tc��IC��L����ܿ���4�P��]|�`   `   �0T���G�E;(��C��o����}�Έ(�#�޾#��<�Y��W+�F�s��F��W+�<�Y�#��#�޾Έ(���}��o���C�E;(���G�`   `   �����iA �k�ɿ�K��~*O�7��<����y��T.�uU��۽ژν�۽uU��T.��y�<���7��~*O��K��k�ɿiA ���`   `   �㿠�ؿ�޼�<!���ye�}M$��X�S)���NK�*x
�sǽf��ӡ��f��sǽ*x
��NK�S)���X�}M$��ye�<!���޼���ؿ`   `   �塿`Y��x�����b�9�/��`�����y��
'�~$߽ܙ���h�KAQ���h�ܙ�}$߽�
'��y�����`�9�/���b�x���`Y��`   `   �Jl�|�c�M���,���	�1�о�U��sES�������wn|��/6�ث��/6�wn|�������sES��U��1�о��	���,�M�|�c�`   `   ��7��2��"���*���M;����>��Q��O����h��<%�=G��<%���h��O���Q���>�M;��*������"��2�`   `   ������������8�Ͼg*���d~���:�	"��`���Hx���5������5��Hx��`��	"���:��d~�g*��8�Ͼ���������`   `   ����T�
	��B�lξ�ݧ��*��[�E�G'��νS����h�,�R��h�S����νG'�[�E��*���ݧ��lξ�B�
	��T�`   `   =�������0^����ھ&�������v�[��,&�%����h½Mǡ��!��Mǡ��h½%����,&�v�[�����&�����ھ0^�������`   `   $)��m%������
�Ӄ�X�ž����<{�n�E����@G�-�轈	߽-��@G����n�E��<{����X�žӃ�
�����m%�`   `   _�7�ů3�dh(�G�Q���AھUj�����>�n��0K�+&5�K�)��&�K�)�+&5��0K�>�n����Uj���AھQ��G�dh(�ů3�`   `   �iD�/P@���4�q�"��8���oǾWۧ�!���4��r�}�;qy�ڂx�;qy�r�}��4��!��Wۧ�oǾ���8�q�"���4�/P@�`   `   M��H��<���*�*��3L ���ܾ[-þ�y���ͱ�q`������lj������q`���ͱ��y��[-þ��ܾ3L �*����*��<��H�`   `   �P�uL�Q@�Q�.�>����cD�S��E徙1� ]���������� ]��1�E�S��cD���>��Q�.�Q@�uL�`   `   �L�`I�<(>�-<.����.�&�k�����U%�>:�!�J�*�P�!�J�>:�U%����k��&�.����-<.�<(>�`I�`   `   C�C��Q@��6��&)�z��mX���č"�o�=���b����K��R��K�������b�o�=�Í"���mX�z���&)��6��Q@�`   `    L5�k\2��v*�X ��h�e.�39%�c�C�T�t�o&���X���6տ$߿�6տ�X��o&��T�t�c�C�39%�e.��h�X ��v*�k\2�`   `   ��"�:t ����{���Y�ϻ���7�n4j�o]���r̿�B ����;������B ��r̿o]��n4j���7�ϻ��Y�{�����:t �`   `   ^��3�	����a�܏ ��[J�'C����w��(�J�G���S�J�G��(�w���'C���[J�܏ �a����	�3�`   `   ѥ��{�oK󾟥��"�Z�=^���_�<��d�P��^|�R���^|�d�P�<���_�=^��Z��"����oK�{���`   `   �žoƾ��ɾ^�־I���G!��Qc�̴���N��_32��bp��S��P����S���bp�_32��N��̴���Qc�G!�I���^�־��ɾoƾ`   `   � ���Ƞ��㧾�C&�dq�&�b�8��LC ���9��^|�Ԛ���٧�Ԛ���^|���9�LC �8��&�b�dq�C&�򺾕㧾�Ƞ�`   `   �z��$�X��-���!.;�����W�,��f���1��<p��P��χ���P���<p��1�f��,����W����!.;-���X���$�`   `   �{?���E�v,[��?��~���Tc��IC��L����ܿ���4�P��]|�m����]|�4�P������ܿ�L���IC�Tc�~����?��v,[���E�`   `   s��F��W+�<�Y�#��#�޾Έ(���}��o���C�E;(���G��0T���G�E;(��C��o����}�Έ(�#�޾#��<�Y��W+�F�`   `   ژν�۽uU��T.��y�<���7��~*O��K��k�ɿiA ��������iA �k�ɿ�K��~*O�7��<����y��T.�uU��۽`   `   ҡ��f��sǽ*x
��NK�S)���X�}M$��ye�<!���޼���ؿ�㿠�ؿ�޼�<!���ye�}M$��X�S)���NK�*x
�sǽf��`   `   KAQ���h�ܙ�}$߽�
'��y�����`�9�/���b�x���`Y���塿`Y��x�����b�9�/��`�����y��
'�}$߽ܙ���h�`   `   ׫��/6�wn|�������sES��U��1�о��	���,�M�|�c��Jl�|�c�M���,���	�1�о�U��sES�������wn|��/6�`   `   �;�	�S�^l����ͽߺ���Q�V܎�T��M�꾛��E!�/�� 4�/��E!���M��T��V܎���Q�ߺ���ͽ^l��	�S�`   `   ��L��?g�Ҭ����߽5� ��$`����
Y¾���p�?!�ǐ-�1�1�ǐ-�?!��p���
Y¾����$`�5� ���߽Ҭ���?g�`   `   ����_�����6��)7���{��K��	�վ�^� }�V�-��F:�f�>��F:�V�-� }��^�	�վ�K����{��)7�6�����_��`   `   ʦ��]�������u&V�G����^������n-��)B���O��eT���O��)B�n-������^��G���u&V������]��`   `   �G齼��V��M�>�,�{�!���9�ؾ35	��<'�"6C���Y�mgh�-wm�mgh���Y�"6C��<'�35	�9�ؾ!���,�{�L�>�V�����`   `   q!��(��?�F�h�ct��n��|��Q;���9�bX��Yp�����˂�����Yp�bX���9�Q;�|��n��ct��F�h��?��(�`   `   �O`�<5f�l_y��ӎ�� �վ~���<'�=�I�Ai��o������ڌ������o��Ai�=�I��<'�~�� �վ��ӎ�l_y�<5f�`   `   �����랾Y���ⰾfȾX�={���1�J|T���t�����t�����t��������t�J|T���1�={�X�fȾ�ⰾY���랾`   `   ��޾gݾi�۾1޾
��ܞ�}���8�L�Y��ly�3ቿ�ϒ�����ϒ�3ቿ�ly�L�Y���8�}�ܞ�
��1޾i�۾gݾ`   `   ӈ�I��� ��4���Bh�^�!�?3;�X@Y���v�����n�������n���������v�X@Y�?3;�^�!�Bh����4�� �I��`   `   �8]�8W���G�Y5��d&��G!�;?(��I:��9S�zm�����ቿ�����ቿ���zm��9S��I:�;?(��G!��d&�Y5���G�8W�`   `   4����C��4\��\�g��H�1�3�:.�-�6�o�H�^���q��B�\���B���q�^�o�H�-�6�:.�1�3��H�\�g�4\���C��`   `   �[̿�ÿM歿�ȑ�C�n�*WH��4� �0��K:�z�I���Y�*e�cDi�*e���Y�z�I��K:� �0��4�*WH�C�n��ȑ�M歿�ÿ`   `   �3��2���`ڿ�����Ћ��-]��9�9�)���)���2��;>��G�hJ��G��;>���2���)�9�)��9��-]��Ћ������`ڿ�2��`   `   �E�,�O7��Ͽ���o�n�t&<�HL!��e�6���'!�_A'�Τ)�_A'��'!�6���e�HL!�t&<�o�n�����ϿO7�,�`   `   ;B4�!�*�����俒����ry��R;��G����^��/��(��	�(�/��^������G��R;��ry����������!�*�`   `   �<���1��+��쿎筿�ay��5�nO�\��2gپ"־��׾��ؾ��׾"־2gپ\��nO��5��ay��筿���+���1�`   `   �F4��{*�>��$�p ���qm�E�(������hɾU����Ԩ��Ħ�ᠦ��Ħ��Ԩ�U����hɾ����E�(��qm�p ���$�>��{*�`   `   r��*�̡��[̿�7���<W���2�۾:����⎾7�����{�b�y���{�7����⎾:���2�۾���<W��7���[̡̿��*�`   `   ��������Iٿ�����:�V������^��mb� VF�F�9�e6�F�9� VF�mb��^�����V����:�����Iٿ����`   `   ��Ͽ}ƿ䭿����:W����W�޾�坾�Qf��2�H���x�2D��x�H���2��Qf��坾W�޾����:W����䭿}ƿ`   `   �����M��+����`�x/����R������`i>��]��߽�O���鷽�O���߽�]�`i>������R����x/���`�+���M��`   `   ��w���n���V��5��R��۾\���Lf��#��l����2u���H��2u������l齖#��Lf�\���۾�R��5���V���n�`   `   ��I�L�C��32�;��$���¾��QpS�(�-нF���d�~N��d�F��-н(�QpS����¾�$��;��32�L�C�`   `   � 4�/��E!���M��T��V܎���Q�ߺ���ͽ^l��	�S��;�	�S�^l����ͽߺ���Q�V܎�T��M�꾛��E!�/�`   `   1�1�ǐ-�?!��p���
Y¾����$`�5� ���߽Ҭ���?g���L��?g�Ҭ����߽5� ��$`����
Y¾���p�?!�ǐ-�`   `   f�>��F:�V�-� }��^�	�վ�K����{��)7�6�����_������_�����6��)7���{��K��	�վ�^� }�V�-��F:�`   `   �eT���O��)B�n-������^��G���u&V������]��ʦ��]�������u&V�G����^������n-��)B���O�`   `   -wm�mgh���Y�"6C��<'�35	�9�ؾ!���,�{�M�>�V������G齼��V��M�>�,�{�!���9�ؾ35	��<'�"6C���Y�mgh�`   `   �˂�����Yp�bX���9�Q;�|��n��ct��F�h��?��(�q!��(��?�F�h�ct��n��|��Q;���9�bX��Yp����`   `   ڌ������o��Ai�=�I��<'�~�� �վ��ӎ�l_y�<5f��O`�<5f�l_y��ӎ�� �վ~���<'�=�I�Ai��o������`   `   ���t��������t�J|T���1�={�X�fȾ�ⰾY���랾�����랾Y���ⰾfȾX�={���1�J|T���t�����t��`   `   ����ϒ�3ቿ�ly�L�Y���8�}�ܞ�
��1޾i�۾gݾ��޾gݾi�۾1޾
��ܞ�}���8�L�Y��ly�3ቿ�ϒ�`   `   ����n���������v�X@Y�?3;�^�!�Bh����4�� �I��ӈ�I��� ��4���Bh�^�!�?3;�X@Y���v�����n���`   `   �����ቿ���zm��9S��I:�;?(��G!��d&�Y5���G�8W��8]�8W���G�Y5��d&��G!�;?(��I:��9S�zm�����ቿ`   `   \���B���q�^�o�H�-�6�:.�1�3��H�\�g�4\���C��4����C��4\��\�g��H�1�3�:.�-�6�o�H�^���q��B�`   `   cDi�*e���Y�z�I��K:�!�0��4�*WH�C�n��ȑ�M歿�ÿ�[̿�ÿM歿�ȑ�C�n�*WH��4� �0��K:�z�I���Y�*e�`   `   hJ��G��;>���2���)�9�)��9��-]��Ћ������`ڿ�2���3��2���`ڿ�����Ћ��-]��9�9�)���)���2��;>��G�`   `   Τ)�_A'��'!�6���e�HL!�t&<�o�n�����ϿO7�,��E�,�O7��Ͽ���o�n�t&<�HL!��e�6���'!�_A'�`   `   �	�(�/��^������G��R;��ry����������!�*�;B4�!�*�����俒����ry��R;��G����^��/��(�`   `   ��ؾ��׾"־2gپ\��nO��5��ay��筿���+���1��<���1��+��쿎筿�ay��5�nO�\��2gپ"־��׾`   `   ᠦ��Ħ��Ԩ�U����hɾ����E�(��qm�p ���$�>��{*��F4��{*�>��$�p ���qm�E�(������hɾU����Ԩ��Ħ�`   `   b�y���{�7����⎾:���2�۾���<W��7���[̡̿��*�r��*�̡��[̿�7���<W���2�۾:����⎾7�����{�`   `   e6�F�9� VF�mb��^�����V����:�����Iٿ������������Iٿ�����:�V������^��mb� VF�F�9�`   `   2D��x�H���2��Qf��坾W�޾����:W����䭿}ƿ��Ͽ}ƿ䭿����:W����W�޾�坾�Qf��2�H���x�`   `   �鷽�O���߽�]�`i>������R����x/���`�+���M�������M��+����`�x/����R������`i>��]��߽�O��`   `   �H��2u������l齖#��Lf�\���۾�R��5���V���n���w���n���V��5��R��۾\���Lf��#��l����2u��`   `   ~N��d�E��-н(�QpS����¾�$��;��32�L�C���I�L�C��32�;��$���¾��QpS�(�-нE���d�`   `   ��u�6{���ұ�[|��O/���q�����jоG�}��T-�f�:���?�f�:��T-�}�G��jо�����q�O/�[|���ұ�6{��`   `   �o��M����KŽ�� G��Ɖ������쾳����+���A�D�O���T�D�O���A���+�����������Ɖ�� G���KŽM���`   `   ���x±��M꽤"%�7�i��P���S׾�3
��)��G�Ӝ_�<@o���t�<@o�Ӝ_��G��)��3
��S׾�P��7�i��"%��M�x±�`   `   ��Ƚ��ݽg��NmE�J뉾�g��V\����!��QF���g��L������(������L����g��QF���!�V\���g��J뉾MmE�g����ݽ`   `   �� �_+��/�uk��L��[�۾���c@:��0c�7��_������	������_���7���0c�c@:����[�۾�L��uk��/�_+�`   `   ��%��f1�T�U����������H���Q$�@�P�Wf}�p���t��7h��H3��7h���t��p��Wf}�@�P��Q$��H����������T�U��f1�`   `   ��U��a��$������5�Ѿ�0
��-4��0c�S��\T��*���Yſ�Y˿Yſ*���\T��S���0c��-4��0
�5�Ѿ�����$���a�`   `   [���Џ��$���׻�.�����Q@�'�o������M������?ӿ�;ڿ�?ӿ����M������'�o�Q@����.�龙׻��$���Џ�`   `   5{��ڐ���Sľb�ھ��4�C�G�W/v�����Ĭ�wYſ�pؿ��߿�pؿwYſ�Ĭ����W/v�C�G�4���b�ھ�Sľڐ��`   `   ��f�y���BP �R,��&�O�J�Z�u�4
�����O���Oӿ�6ڿ�Oӿ�O����4
��Z�u�O�J��&�R,�BP �y����f�`   `   ���C��z����N
��U-�V�I��Bo�!c��[���+���Zſ�2˿Zſ+���[���!c���Bo�V�I��U-�N
�����z��C�`   `   �O��K��@��4��.�HS3�3�E��uc�@Q��OY��(祿��������(祿OY��@Q���uc�2�E�HS3��.��4��@��K�`   `   �9��FY���l�hT���@��9�+�?���S��Do��Z�������眿iV���眿�����Z���Do���S�+�?��9���@�hT��l�FY��`   `   O|������Í�(�u���S�}>�1#8��A�?T�b-k�D��H_��W ��H_��D��b-k�?T��A�1#8�}>���S�(�u��Í����`   `   �C��R���/����"�c���@��/��Z-�]�7���G��W��6c�E_g��6c��W���G�]�7��Z-��/���@�"�c����/�R���`   `   �!ҿ�7ɿ�±�ځ����l���?�?n$�hx�7<�C^$��j/�T�7�;�T�7��j/�C^$�6<�hx�?n$���?���l�ځ���±��7ɿ`   `   �]ٿe�Ͽ���� ���l���9���������
��9
���������9
��
����������9��l�� �����e�Ͽ`   `   �3ҿ��ȿA������b�a���-��'	���̩Ӿ
)оuԾ�پ�;ܾ�پuԾ
)о̩Ӿ���'	���-�b�a����A�����ȿ`   `   J߾��������9��reN�I��s�fľ۫��p�������\���0���\�����p���۫��fľ�s�I�reN��9��������`   `   @���m���"����g���5��
�óҾ|��������y���m�nj�	�i�nj���m��y�����|���óҾ�
���5���g�"��m���`   `   �����h����l�UF�G��"������K���>a�[s@��"/�]['��6%�]['��"/�[s@��>a��K�������"�G�UF���l��h��`   `   �e�I�]�	'H���)�	��Ծ�l���dt�$�<������P��C��P�ｧ����$�<��dt��l���Ծ	���)�	'H�I�]�`   `   ��F�}�@�l�/�T��U-���_ľ���>8a�Q�(�q� ��Kνa౽#֨�a౽�Kνq� �Q�(�>8a�����_ľU-��T��l�/�}�@�`   `   �T:�[85�%�&����C{󾬮¾8��Ym`�-`$����������������������-`$�Ym`�8����¾C{���%�&�[85�`   `   ��?�f�:��T-�}�G��jо�����q�O/�[|���ұ�6{����u�6{���ұ�[|��O/���q�����jоG�}��T-�f�:�`   `   ��T�D�O���A���+�����������Ɖ�� G���KŽM����o��M����KŽ�� G��Ɖ������쾳����+���A�D�O�`   `   ��t�<@o�Ӝ_��G��)��3
��S׾�P��7�i��"%��M�x±����x±��M꽤"%�7�i��P���S׾�3
��)��G�Ӝ_�<@o�`   `   �(������L����g��QF���!�V\���g��J뉾NmE�g����ݽ��Ƚ��ݽg��NmE�J뉾�g��V\����!��QF���g��L�����`   `   	������_���7���0c�c@:����[�۾�L��uk��/�_+��� �_+��/�uk��L��[�۾���c@:��0c�7��_������`   `   H3��8h���t��p��Wf}�@�P��Q$��H����������T�U��f1���%��f1�T�U����������H���Q$�@�P�Wf}�p���t��7h��`   `   �Y˿Yſ*���\T��S���0c��-4��0
�5�Ѿ�����$���a���U��a��$������5�Ѿ�0
��-4��0c�S��\T��*���Yſ`   `   �;ڿ�?ӿ����M������'�o�Q@����.�龙׻��$���Џ�[���Џ��$���׻�.�����Q@�'�o������M������?ӿ`   `   ��߿�pؿwYſ�Ĭ����W/v�C�G�4���b�ھ�Sľڐ��5{��ڐ���Sľb�ھ��4�C�G�W/v�����Ĭ�wYſ�pؿ`   `   �6ڿ�Oӿ�O����4
��Z�u�O�J��&�R,�BP �y����f��f�y���BP �R,��&�O�J�Z�u�4
�����O���Oӿ`   `   �2˿Zſ+���[���!c���Bo�V�I��U-�N
�����z��C����C��z����N
��U-�V�I��Bo�!c��[���+���Zſ`   `   ������(祿OY��@Q���uc�3�E�HS3��.��4��@��K��O��K��@��4��.�HS3�3�E��uc�@Q��OY��(祿��`   `   iV���眿�����Z���Do���S�+�?��9���@�hT��l�FY���9��FY���l�hT���@��9�+�?���S��Do��Z�������眿`   `   W ��H_��D��b-k�?T��A�1#8�}>���S�(�u��Í����O|������Í�(�u���S�}>�1#8��A�?T�b-k�D��H_��`   `   E_g��6c��W���G�]�7��Z-��/���@�"�c����/�R����C��R���/����"�c���@��/��Z-�]�7���G��W��6c�`   `   ;�T�7��j/�C^$�7<�hx�?n$���?���l�ځ���±��7ɿ�!ҿ�7ɿ�±�ځ����l���?�?n$�hx�7<�C^$��j/�T�7�`   `   ������9
��
����������9��l�� �����e�Ͽ�]ٿe�Ͽ���� ���l���9���������
��9
���`   `   �;ܾ�پuԾ
)о̩Ӿ���'	���-�b�a����A�����ȿ�3ҿ��ȿA������b�a���-��'	���̩Ӿ
)оuԾ�پ`   `   �0���\�����p���۫��fľ�s�I�reN��9��������J߾��������9��reN�I��s�fľ۫��p�������\��`   `   	�i�nj���m��y�����|���óҾ�
���5���g�"��m���@���m���"����g���5��
�óҾ|��������y���m�nj�`   `   �6%�]['��"/�[s@��>a��K�������"�G�UF���l��h�������h����l�UF�G��"������K���>a�[s@��"/�]['�`   `   C��P�ｧ����$�<��dt��l���Ծ	���)�	'H�I�]��e�I�]�	'H���)�	��Ծ�l���dt�$�<������P��`   `   #֨�a౽�Kνq� �Q�(�>8a�����_ľU-��T��l�/�}�@���F�}�@�l�/�T��U-���_ľ���>8a�Q�(�q� ��Kνa౽`   `   ������������-`$�Ym`�8����¾C{���%�&�[85��T:�[85�%�&����C{󾬮¾8��Ym`�-`$����������`   `   %s��!!��w�ܽJ�$pQ�T㎾:w����O�0��GF�dU��(Z�dU��GF�0��O���:w��T㎾$pQ�J�w�ܽ!!��`   `   m8��<���F��,�-���u��詾7(�����3��fS�k�l���}�¿����}�k�l��fS���3���7(��詾��u�,�-�F��<���`   `   7GŽݽܽ����N�=𒾇4̾N	�)�0�]�X�Ry}�᥍�ۜ��V(��ۜ��᥍�Ry}�]�X�)�0�N	��4̾=𒾬�N���ݽܽ`   `   *j�����X/�
tv�&Ǯ�V��e#���Q�������߀�����%�����߀����������Q��e#�V�&Ǯ�
tv��X/����`   `   &c�4�"�6]Q�����/̾����=��gr��˓����O�ȿ��ܿ�{���ܿO�ȿ����˓��gr���=����/̾���6]Q�4�"�`   `   ��3�yD���v�Mg������ �%�U�Kԇ��æ�=uɿ4��̦�OZ�̦�4��=uɿ�æ�Kԇ�%�U�� ����Mg����v�yD�`   `   ��Y�N|j��L���j���r�ʓ0��Hi��˓�Ɵ���C�0�	�����$���0�	��C�Ɵ���˓��Hi�ʓ0��r��j���L��N|j�`   `   ����������Ҿ�t���<�3�v�c
����ÿܵ�������.��J7���.����ܵ����ÿb
��3�v���<��t��Ҿ�����`   `   �Ο�릾�����羳J�
%D��w}�:���ڦȿy:��C�5��>>�5�C�y:��ڦȿ:����w}�
%D��J�������릾`   `   4$þ��Ⱦ�oھ���f8�0G�@}����ĿXl�����.��F7��.���Xl����Ŀ�@}�0G�f8�����oھ��Ⱦ`   `   7ﾉ��4���ζ
�}�!��FF�I�v�����eɹ�/}俄�	�c��i$�c���	�/}�eɹ�����I�v��FF�}�!�ζ
�4������`   `   8������z�	����&��;B�A~j�}���<ө��ʿ}R�j}�y�j}�}R��ʿ<ө�}���A~j��;B���&�	���z����`   `   g�/��z-�a�(�� &�7�*���;��+Z����מ���'��x�ȿ��ۿ�E㿰�ۿx�ȿ�'��מ������+Z���;�7�*�� &�a�(��z-�`   `   � N�1�I��?���3�vW.��4�qG�e�m���ɖ�s���]*���Ӹ�]*��s����ɖ�m��e�qG��4�vW.���3��?�1�I�`   `   �h���b�ՀR�?���/���*�/�2�}LF�*a�)}��,��Iϓ� Iϓ��,��)}�*a�}LF�/�2���*���/�?�ՀR���b�`   `   Ql{���s�|B_�MuE��l.�Oe ��Z���'���9��N���a���n��s���n���a��N���9���'��Z�Oe ��l.�MuE�|B_���s�`   `   ���Kny�̘b��D���(�WU�K�
�	���T��#�(�0�e]:���=�e]:�(�0��#��T�	��K�
�WU���(��D�̘b�Kny�`   `   �{�G�r���[�Q!=����6��m�����������[��zG�[�����������m��6�����Q!=���[�G�r�`   `   ��j�ߖb�!�L��/������ҾϾ����*2��5����gžcC̾e�ξcC̾�gž5���*2������ҾϾ������/�!�L�ߖb�`   `   �IT��=M��:�*���K�Nؾ��� ��B�������E䏾M8��+E��M8��E䏾����B���� ����Nؾ�K�*���:��=M�`   `   q?��9��(����N�փľY���_���)�j�AY���Q��-O���N��-O���Q�AY�)�j�_���Y���փľN����(��9�`   `   �;1��,����Ʀ	��澚����O���p�|G�p�+�T��N����N��T��p�+�|G��p��O��������Ʀ	�����,�`   `   �/���*�����
�w��b����(���j���7��~�@d����ܽ�mԽ��ܽ@d���~���7��j��(��b���w���
������*�`   `   �=��f8��+��I�����о�|����y���;��_�W۽�/��},���/��W۽�_���;���y��|���о����I��+��f8�`   `   �(Z�dU��GF�0��O���:w��T㎾$pQ�K�w�ܽ!!��%s��!!��w�ܽK�$pQ�T㎾:w����O�0��GF�dU�`   `   ¿����}�k�l��fS���3���7(��詾��u�,�-�F��<���m8��<���F��,�-���u��詾7(�����3��fS�k�l���}�`   `   V(��ۜ��᥍�Ry}�]�X�)�0�N	��4̾=𒾬�N���ݽܽ7GŽݽܽ����N�=𒾇4̾N	�)�0�]�X�Ry}�᥍�ۜ��`   `   %�����߀����������Q��e#�V�&Ǯ�
tv��X/����*j�����X/�
tv�&Ǯ�V��e#���Q�������߀�����`   `   �{���ܿO�ȿ����˓��gr���=����/̾���6]Q�4�"�&c�4�"�6]Q�����/̾����=��gr��˓����O�ȿ��ܿ`   `   OZ�̦�4��=uɿ�æ�Kԇ�%�U�� ����Mg����v�yD���3�yD���v�Mg������ �%�U�Kԇ��æ�=uɿ4��̦�`   `   ��$���0�	��C�Ɵ���˓��Hi�ʓ0��r��j���L��N|j���Y�N|j��L���j���r�ʓ0��Hi��˓�Ɵ���C�0�	���`   `   �J7���.����ܵ����ÿc
��3�v���<��t��Ҿ���������������Ҿ�t���<�3�v�c
����ÿܵ�������.�`   `   �>>�5�C�y:��ڦȿ:����w}�
%D��J�������릾�Ο�릾�����羳J�
%D��w}�:���ڦȿy:��C�5�`   `   �F7��.���Xl����Ŀ�@}�0G�f8�����oھ��Ⱦ4$þ��Ⱦ�oھ���f8�0G�@}����ĿXl�����.�`   `   �i$�c���	�/}�eɹ�����I�v��FF�}�!�ζ
�4������7ﾉ��4���ζ
�}�!��FF�I�v�����eɹ�/}俄�	�c�`   `   y�j}�}R��ʿ<ө�}���A~j��;B���&�	���z����8������z�	����&��;B�A~j�}���<ө��ʿ}R�j}�`   `   �E㿰�ۿx�ȿ�'��מ������+Z���;�7�*�� &�a�(��z-�g�/��z-�a�(�� &�7�*���;��+Z����מ���'��x�ȿ��ۿ`   `   �Ӹ�]*��s����ɖ�m��e�qG��4�vW.���3��?�1�I�� N�1�I��?���3�vW.��4�qG�e�m���ɖ�s���]*��`   `    Iϓ��,��)}�*a�}LF�/�2���*���/�?�ՀR���b��h���b�ՀR�?���/���*�/�2�}LF�*a�)}��,��Iϓ�`   `   �s���n���a��N���9���'��Z�Oe ��l.�MuE�|B_���s�Ql{���s�|B_�MuE��l.�Oe ��Z���'���9��N���a���n�`   `   ��=�e]:�(�0��#��T�	��K�
�WU���(��D�̘b�Kny����Kny�̘b��D���(�WU�K�
�	���T��#�(�0�e]:�`   `   zG�[�����������m��6�����Q!=���[�G�r��{�G�r���[�Q!=����6��m�����������[��`   `   e�ξcC̾�gž5���*2������ҾϾ������/�!�L�ߖb���j�ߖb�!�L��/������ҾϾ����*2��5����gžcC̾`   `   +E��M8��E䏾����B���� ����Nؾ�K�*���:��=M��IT��=M��:�*���K�Nؾ��� ��B�������E䏾M8��`   `   ��N��-O���Q�AY�)�j�_���Y���փľN����(��9�q?��9��(����N�փľY���_���)�j�AY���Q��-O�`   `   ��M��T��p�+�|G��p��O��������Ʀ	�����,��;1��,����Ʀ	��澚����O���p�|G�p�+�T��M��`   `   �mԽ��ܽ@d���~���7��j��(��b���w���
������*��/���*�����
�w��b����(���j���7��~�@d����ܽ`   `   },���/��W۽�_���;���y��|���о����I��+��f8��=��f8��+��I�����о�|����y���;��_�W۽�/��`   `   ��½Q�Խ���
5�|�x�+��U�߾13���/���N���g�4?x���}�4?x���g���N���/�13�U�߾+��|�x�
5����Q�Խ`   `   ��ν�)�j��^�R������]ξ�e
�O:2���Z����?E��%z��_��%z��?E�������Z�O:2��e
��]ξ����^�R�i���)�`   `   �;�u���w1�q|��#��B�����)�G�Z�Y��������O���|��v.ƿ�|���O������Y���G�Z���)�B����#��q|��w1�u��`   `   ��s��VYS��7���r׾�1��K�ZC��M蟿�῿���m���!S�m�����࿽῿M蟿ZC���K��1��r׾�7��VYS�s��`   `   �p*�!�=���x�
꯾����0�"�l��&��Ĵ������i��&�j4/��&��i����Ĵ���&��"�l��0����	꯾��x�!�=�`   `   ��H�&^�A���
ɾ�0���G�턿�u��_�޿���9�M�X���d�M�X��9���_�޿�u��턿��G��0�
ɾA���&^�`   `   ��h�w\��`����߾���"�Z�hܐ�:�������f.��a�qS��̋�qS���a��f.����9���hܐ�"�Z������߾�`��w\�`   `   u������g�������)���g�'���
˿΄�c(C���}�~���f+��~�����}�c(C�΄��
˿'����g��)����g�������`   `   Sȗ�����4�ľ� ���/�b)n�/����oпj�WK��S�����Zܤ�����S��WK�j��oп/���b)n���/�� �4�ľ����`   `   *@��>뵾��Ծ���g�2�/n�X,��7�̿��C�TG~�����#'������TG~��C��7�̿X,��/n�g�2������Ծ>뵾`   `   D�þ�q˾!��j�
�ݧ1���g����}�����4/��a�kS��A���kS���a��4/���}�������g�ݧ1�j�
�!���q˾`   `   a�ݾ�I���������-��E\��a��{l����῱n���9�A{X�d�A{X���9��n����{l���a���E\��-���������I�`   `   �������*��L�x�'�_�L�`�}��2��s~��o���j�,Z&�g.�,Z&��j�o��s~���2��`�}�_�L�x�'�L�*�����`   `   ��
���
����,p����M�:�xa��E������$�����߿���<������߿$��������E��xa�M�:����,p������
�`   `   �J�������j�U�|�'��:C�1�g�k3��e��� ���P���d	ÿP��� ���e���k3��1�g��:C�|�'�U��j������`   `   G�Ӌ��e�hW������ͤ%���?�y�^��A}�����������������A}�y�^���?�ͤ%������hW��e�Ӌ�`   `   s� ��k�,����
����� �G�
������/�D�F���Z���g���l���g���Z�D�F���/����G�
�� ������
�,���k�`   `   �`�������m?��k�-��y羋i��^��h��|$��.�A{1��.�|$�h��^���i���y�-澾k�m?�������`   `   ���D����
������!߾&�˾z¾��ľn�Ͼ�߾*'����, ���*'��߾n�Ͼ��ľz¾&�˾�!߾������
�D��`   `   ��E�����@�о� ��$���m����:��x���r�������WŴ�����r���x����:��m���$���� ��@�о�����E�`   `   Ei�a�����+��E}˾t����ٗ��V������y� y�{�*-|�{� y��y�����V���ٗ�t���E}˾+�꾆��a��`   `   �D����]
���+�Ӿ���������9{�:/Z���D�w�8�a�2��(1�a�2�w�8���D�:/Z��9{���������+�Ӿ��]
����`   `   U�+��'�e��Ҽ
��X�r�ľ�A��<�'5N�Q�*�N���u����N�Q�*�'5N�<��A��r�ľ�X�Ҽ
�e���'�`   `   ��M�;I��P;�]�&�k���|�IG��jx��^XY�(v&�H��J�޽NyѽJ�޽H��(v&�^XY�jx��IG���|�k��]�&��P;�;I�`   `   ��}�4?x���g���N���/�13�U�߾+��|�x�
5����Q�Խ��½Q�Խ���
5�|�x�+��U�߾13���/���N���g�4?x�`   `   _��%z��?E�������Z�O:2��e
��]ξ����^�R�j���)���ν�)�j��^�R������]ξ�e
�O:2���Z����?E��%z��`   `   v.ƿ�|���O������Y���G�Z���)�B����#��q|��w1�u���;�u���w1�q|��#��B�����)�G�Z�Y��������O���|��`   `   !S�m�����࿽῿M蟿ZC���K��1��r׾�7��VYS�s����s��VYS��7���r׾�1��K�ZC��M蟿�῿���m���`   `   j4/��&��i����Ĵ���&��"�l��0����
꯾��x�!�=��p*�!�=���x�
꯾����0�"�l��&��Ĵ������i��&�`   `   ��d�M�X��9���_�޿�u��턿��G��0�
ɾA���&^���H�&^�A���
ɾ�0���G�턿�u��_�޿���9�M�X�`   `   ̋�qS���a��f.����:���hܐ�"�Z������߾�`��w\���h�w\��`����߾���"�Z�hܐ�:�������f.��a�qS��`   `   f+��~�����}�c(C�΄��
˿'����g��)����g�������u������g�������)���g�'���
˿΄�c(C���}�~���`   `   Zܤ�����S��WK�j��oп/���b)n���/�� �4�ľ����Sȗ�����4�ľ� ���/�b)n�/����oпj�WK��S�����`   `   #'������TG~��C��7�̿X,��/n�g�2������Ծ>뵾*@��>뵾��Ծ���g�2�/n�X,��7�̿��C�TG~�����`   `   A���kS���a��4/���}�������g�ݧ1�j�
�!���q˾D�þ�q˾!��j�
�ݧ1���g����}�����4/��a�kS��`   `   d�A{X���9��n����{l���a���E\��-���������I�a�ݾ�I���������-��E\��a��{l����῱n���9�A{X�`   `   g.�,Z&��j�o��s~���2��`�}�_�L�x�'�L�*������������*��L�x�'�_�L�`�}��2��s~��o���j�,Z&�`   `   <������߿$��������E��xa�M�:����,p������
���
���
����,p����M�:�xa��E������$�����߿���`   `   d	ÿP��� ���e���k3��1�g��:C�|�'�U��j�������J�������j�U�|�'��:C�1�g�k3��e��� ���P���`   `   ����������A}�y�^���?�ͤ%������hW��e�Ӌ�G�Ӌ��e�hW������ͤ%���?�y�^��A}�������`   `   ��l���g���Z�D�F���/����G�
�� ������
�,���k�s� ��k�,����
����� �G�
������/�D�F���Z���g�`   `   A{1��.�|$�h��^���i���y�-澾k�m?��������`�������m?��k�-��y羋i��^��h��|$��.�`   `   �, ���+'��߾n�Ͼ��ľz¾&�˾�!߾������
�D�����D����
������!߾&�˾z¾��ľn�Ͼ�߾+'���`   `   WŴ�����r���x����:��m���$���� ��@�о�����E���E�����@�о� ��$���m����:��x���r�������`   `   *-|�{� y��y�����V���ٗ�t���E}˾+�꾆��a��Ei�a�����+��E}˾t����ٗ��V������y� y�{�`   `   �(1�a�2�w�8���D�:/Z��9{���������+�Ӿ��]
�����D����]
���+�Ӿ���������9{�:/Z���D�w�8�a�2�`   `   t����N�Q�*�'5N�<��A��r�ľ�X�Ҽ
�e���'�U�+��'�e��Ҽ
��X�r�ľ�A��<�'5N�Q�*�N���`   `   NyѽJ�޽H��(v&�^XY�jx��IG���|�k��]�&��P;�;I���M�;I��P;�]�&�k���|�IG��jx��^XY�(v&�H��J�޽`   `   ����p��M@�SMS�[͐�Y�ľ�h�� '�P�L���o�����e��ɲ���e�������o�P�L�� '��h�Y�ľ[͐�SMS�M@��p��`   `   7������1�+�w��K��֬�C�#���R�D�������a��a��쒽�a���a�����D�����R�C�#�֬�K��+�w��1���`   `   _�4�w�P�����n�վ��TpJ�R���;W���T����߿�������������߿�T��;W��R���TpJ���n�վ����w�P�4�`   `   ��%���9�ow��I���. �K�4�2�r�����Lſė�����c�2��$<�c�2����ė���Lſ���2�r�J�4��. ��I��ow���9�`   `   b�B��Z�s�PSϾ�
���R��܌�p~���f���'���W���}������}���W��'��f��p~���܌���R��
�OSϾs��Z�`   `   �Sa�1'{����'��>F*�2�m��7��5ؿ�0�>Z�6/���M������M��6/��>Z��0�5ؿ�7��2�m�>F*�'�����1'{�`   `   ��~��S���[���a���:�飁��2���e��\�8�w���:D��A�������A���:D��w���\�8��e���2��飁���:��a��[���S��`   `   �?��2����Ⱦ���&�F�M���*���ڎ��?O�6=������/������/������6=���?O�ڎ�)���M���&�F�����Ⱦ2���`   `   Sə�"秾�Ծؿ�a�L�*6��zR���:���W�fٝ�;���0��
�0��;���fٝ���W��:�zR��*6��a�L�ؿ��Ծ"秾`   `   RU�������yܾR�E�L�l#��X8��%@���O��������N@�����N@�����������O�%@�X8��l#��E�L�R��yܾ����`   `   �K��",������)�z�G�v��`E��������9����`���Մ���X��Մ��`��������9�����`E��u��z�G��)����",��`   `   @⺾��ľs����t=��{�����qۿ.��C[��b��;��<���;���b��C[�.��qۿ�����{��t=���s���ľ`   `   
�ľ��̾@]�)
���/���d����?��)���IS(�i�W��}�t����}�i�W�IS(�)���?�������d���/�)
�@]征�̾`   `   )�;`$Ӿ��;~��k ���J��\��CΟ��ǿ�P��^����1�f�:���1�^���P���ǿCΟ��\����J��k �;~���`$Ӿ`   `   ��ԾȰ׾��᾿A���O���/���Z��	���+��,W���}޿1j���� �1j���}޿,W���+���	����Z���/��O��A�����Ȱ׾`   `   I�ؾ	�پ��ݾh�辐� �X�R5�vY[�� ��S
��e᧿�紿�����紿e᧿S
��� ��vY[�R5�X��� �h�辛�ݾ	�پ`   `   	ھپ:�׾ھ�d復���1��6.�
�L��j�����e�㌿e󉿀����j�
�L��6.��1�����d�ھ:�׾پ`   `   ��پ�Z׾U�Ѿ>;9�;/Aؾ�V�����T�2j1�X�C�?�O�_�S�?�O�X�C�2j1��T�����V�/Aؾ9�;>;U�Ѿ�Z׾`   `   ��ھ�׾�7Ͼ��ľ`��9:��3�þ�2Ծq@��n�����8�������n�q@��2Ծ3�þ9:��`����ľ�7Ͼ�׾`   `   6㾢�޾@�Ӿ��ľ�Y������2s���1��B�������t}ʾ�4ӾHe־�4Ӿt}ʾ����B����1��2s�������Y����ľ@�Ӿ��޾`   `   pB��A��b徍�Ѿd8��B���"ܙ��ߐ��i��l���ؐ�����䀹������ؐ�l���i���ߐ�"ܙ�B���d8����Ѿ�b�A�`   `   ��.����h��Ҿ�h��a���/w���'r��`�q$V�֤Q�2iP�֤Q�q$V��`��'r�/w��a����h���Ҿ�h��.��`   `   �4�+�/��c$�v/�����,Ծ�ۭ��d���g��C��*��L�=���L��*��C��g��d���ۭ��,Ծ���v/��c$�+�/�`   `   Jf�w�`�mR�lz;��' ��z���о����x�A@�Ő��7������7�Ő�A@��x������о�z��' �lz;�mR�w�`�`   `   ɲ���e�������o�P�L�� '��h�Y�ľ[͐�SMS�N@��p������p��N@�SMS�[͐�Y�ľ�h�� '�P�L���o�����e��`   `   쒽�a���a�����D�����R�B�#�֬�K��+�w��1���7������1�+�w��K��֬�B�#���R�D�������a��a��`   `   ���������߿�T��;W��R���TpJ���n�վ����w�P�4�_�4�w�P�����n�վ��TpJ�R���;W���T����߿����`   `   �$<�c�2����ė���Lſ���2�r�J�4��. ��I��ow���9���%���9�ow��I���. �J�4�2�r�����Lſė�����c�2�`   `   �����}���W��'��f��p~���܌���R��
�PSϾs��Z�b�B��Z�s�PSϾ�
���R��܌�p~���f���'���W���}�`   `   ����M��6/��>Z��0�5ؿ�7��2�m�>F*�'�����1'{��Sa�1'{����'��>F*�2�m��7��5ؿ�0�>Z�6/���M��`   `   ����A���:D��w���\�8��e���2��飁���:��a��[���S����~��S���[���a���:�飁��2���e��\�8�w���:D��A���`   `   ����/������6=���?O�ڎ�)���M���&�F�����Ⱦ2����?��2����Ⱦ���&�F�M���)���ڎ��?O�6=������/��`   `   
�0��;���fٝ���W��:�zR��*6��a�L�ؿ��Ծ"秾Sə�"秾�Ծؿ�a�L�*6��zR���:���W�fٝ�;���0��`   `   ���N@�����������O�%@�X8��l#��E�L�R��yܾ����RU�������yܾR�E�L�l#��X8��%@���O��������N@��`   `   �X��Մ��`��������9�����`E��v��z�G��)����",���K��",������)�z�G�v��`E��������9����`���Մ��`   `   <���;���b��C[�.��qۿ�����{��t=���s���ľ@⺾��ľs����t=��{�����qۿ.��C[��b��;��`   `   t����}�i�W�IS(�)���?�������d���/�)
�@]征�̾
�ľ��̾@]�)
���/���d����?��)���IS(�i�W��}�`   `   f�:���1�^���P���ǿCΟ��\����J��k �;~���`$Ӿ)�;`$Ӿ��;~��k ���J��\��CΟ��ǿ�P��^����1�`   `   �� �1j���}޿,W���+���	����Z���/��O��A�����Ȱ׾��ԾȰ׾��᾿A���O���/���Z��	���+��,W���}޿1j��`   `   �����紿e᧿S
��� ��vY[�R5�X��� �h�辛�ݾ	�پI�ؾ	�پ��ݾh�辐� �X�R5�vY[�� ��S
��e᧿�紿`   `   ㌿e󉿀����j�
�L��6.��1�����d�ھ:�׾پ	ھپ:�׾ھ�d復���1��6.�
�L��j�����e�`   `   _�S�?�O�X�C�2j1��T�����V�/Aؾ9�;>;U�Ѿ�Z׾��پ�Z׾U�Ѿ>;9�;/Aؾ�V�����T�2j1�X�C�?�O�`   `   8�������n�q@��2Ծ3�þ9:��`����ľ�7Ͼ�׾��ھ�׾�7Ͼ��ľ`��9:��3�þ�2Ծq@��n�����`   `   He־�4Ӿt}ʾ����B����1��2s�������Y����ľ@�Ӿ��޾6㾢�޾@�Ӿ��ľ�Y������2s���1��B�������t}ʾ�4Ӿ`   `   䀹������ؐ�l���i���ߐ�"ܙ�B���d8����Ѿ�b�A�pB��A��b徍�Ѿd8��B���"ܙ��ߐ��i��l���ؐ�����`   `   2iP�֤Q�q$V��`��'r�/w��a����h���Ҿ�h��.����.����h��Ҿ�h��a���/w���'r��`�q$V�֤Q�`   `   =���L��*��C��g��d���ۭ��,Ծ���v/��c$�+�/��4�+�/��c$�v/�����,Ծ�ۭ��d���g��C��*��L�`   `   �����7�Ő�A@��x������о�z��' �lz;�mR�w�`�Jf�w�`�mR�lz;��' ��z���о����x�A@�Ő��7�`   `   d!�X����1��@n�K=���(޾����=�qGg����J8���V���\���V��J8�����qGg��=�����(޾K=���@n���1�X��`   `   ��
����yH��J����ƾ
�
���:�c�o�����O���:�ǿ��ۿ�g㿂�ۿ:�ǿO�������c�o���:�
�
���ƾ�J���yH���`   `   ����1��l�ǵ��Iw�t�+���f�4哿����ݣ�5:���!�Z�)���!�5:�ݣ翽���4哿��f�t�+�Iw�Ƶ���l��1�`   `   +:�Q�9Ջ���ɾ����N��N��|񴿧���"��[Q�N�u��܁�N�u��[Q���"����|��N���N������ɾ9Ջ�Q�`   `   lY�{t�2���뾃�+�Gop��ס��:޿I� ��e�4���F_������F_��4����e�I� ��:޿�ס�Gop���+���2��{t�`   `   � y�Np��6ѹ����@^B�Rl���׹����/�P�瑘�����o������o�������瑘�/�P�����׹�Rl��@^B����6ѹ�Np��`   `   ����=��V�;(��p�T��⓿�@пq� �/�~��!������&����&�������!��/�~�q� ��@п�⓿p�T�(��V�;�=��`   `   �c���?����ܾ�j�{a��u������E3��e���v����z�%�ۊ.�z�%����v���e���E3�����u��{a��j���ܾ�?��`   `   Sڠ��±�ʷ���"��?g����j���l:�����q������>,���5��>,���q��������l:�j������?g���"�ʷ澆±�`   `   {h��&���3��#�R�e�!��}Q�!�3��Ɛ�^�������%�߆.��%����^����Ɛ�!�3�}Q�!��R�e�#�3��&���`   `   �V���P���`�Y���]��4��k�ҿ4�!�v������>�����������>������v��4�!�k�ҿ�4����]�Y��`��P��`   `   l���6�����oV�&�O�[��w���D	��Q�*���*������'�������*��*���Q��D	�w��[��&�O�oV���㾙6��`   `   ������v�ھ���'[=��Z}��Z���k�+�!��e�/��������!������/����e�+�!��k��Z���Z}�'[=����v�ھ���`   `   �����T��˭Ͼ$� ��P(��+^�؎���D��&s��@#�,Q�i�t�8��i�t�,Q��@#�&s�D��؎���+^��P(�$� �˭Ͼ�T��`   `   ���Dد���þ��龧��^=��`r��8��������g��� ��[(�� �g���翥����8���`r�^=���������þDد�`   `   J��Id��ٸ�ɻҾ�2��v���F���u�or��ج�(�ſ(�ؿ�$�(�ؿ(�ſج�or����u��F�v���2��ɻҾٸ�Id��`   `   [��DL���ٯ��x����ھ2K�d�"B��Kg�@%���铿Z&��3ޡ�Z&���铿@%���Kg�"B�c�1K���ھ�x���ٯ�DL��`   `   [.������,��J���M����ؾK�����P�/���I���^�l�l�c�q�l�l���^���I�P�/���K�����ؾ�M��J��,������`   `   �˰��ٯ�jۭ����
[���^���̾X���A�
��.�!�Ù+�A/�Ù+�.�!�
���A�X���̾�^��
[�����jۭ��ٯ�`   `   �ľ�:¾+������_]��ŵ��g⭾'A��M�ž�־F��k�𾽎��k��F���־M�ž'A��g⭾ŵ��_]�����+����:¾`   `   %��k�徍�ھ�&˾�]��׀��D�����S��~����I���A���ɨ��A���I��~����S������D׀���]���&˾��ھk��`   `   ���҇�6�{��O�ھ;¾���3���o���gy���p���l��k���l���p��gy�o��3�����;¾�O�ھ{��6�҇�`   `   o�A�m_=�.D1�'��	�+��佾O��H���Y���?���1�P-���1���?��Y�H��O��佾+���	�'�.D1�m_=�`   `   ��~��0y��(i���P�~�2�
��	�@˴�����W��-����i������-��W����@˴�	�
��~�2���P��(i��0y�`   `   �\���V��I8�����qGg��=�����(޾K=���@n���1�X��d!�X����1��@n�K=���(޾����=�qGg����I8���V��`   `   �g㿂�ۿ:�ǿO�������c�o���:�
�
���ƾ�J���yH�����
����yH��J����ƾ
�
���:�c�o�����O���:�ǿ��ۿ`   `   Z�)���!�5:�ݣ翽���4哿��f�t�+�Iw�ǵ���l��1�����1��l�ǵ��Iw�t�+���f�4哿����ݣ�5:���!�`   `   �܁�N�u��[Q���"����|��N���N������ɾ9Ջ�Q�+:�Q�9Ջ���ɾ����N��N��|񴿧���"��[Q�N�u�`   `   ����F_��4����e�I� ��:޿�ס�Gop���+���2��{t�lY�{t�2���뾃�+�Gop��ס��:޿I� ��e�4���F_��`   `   ���o�������瑘�/�P�����׹�Rl��@^B����6ѹ�Np��� y�Np��6ѹ����@^B�Rl���׹����/�P�瑘�����o���`   `   ��&�������!��/�~�q� ��@п�⓿p�T�(��V�;�=������=��V�;(��p�T��⓿�@пq� �/�~��!������&��`   `   ۊ.�z�%����v���e���E3�����u��{a��j���ܾ�?���c���?����ܾ�j�{a��u������E3��e���v����z�%�`   `   ��5��>,���q��������l:�j������?g���"�ʷ澆±�Sڠ��±�ʷ���"��?g����j���l:�����q������>,�`   `   ߆.��%����^����Ɛ�!�3�}Q�!��R�e�#�3��&���{h��&���3��#�R�e�!��}Q�!�3��Ɛ�^�������%�`   `   ������>������v��4�!�k�ҿ�4����]�Y��`��P���V���P���`�Y���]��4��k�ҿ4�!�v������>�����`   `   '�������*��*���Q��D	�w��[��&�O�oV���㾙6��l���6�����oV�&�O�[��w���D	��Q�*���*������`   `   �!������/����e�+�!��k��Z���Z}�'[=����v�ھ���������v�ھ���'[=��Z}��Z���k�+�!��e�/�������`   `   8��i�t�-Q��@#�&s�D��؎���+^��P(�%� �˭Ͼ�T�������T��˭Ͼ%� ��P(��+^�؎���D��&s��@#�-Q�i�t�`   `   �[(�� �g���翥����8���`r�^=���������þDد����Dد���þ��龧��^=��`r��8��������g��� �`   `   �$�(�ؿ(�ſج�or����u��F�v���2��ɻҾٸ�Id��J��Id��ٸ�ɻҾ�2��v���F���u�or��ج�(�ſ(�ؿ`   `   4ޡ�Z&���铿@%���Kg�"B�d�2K���ھ�x���ٯ�DL��[��DL���ٯ��x����ھ2K�d�"B��Kg�@%���铿Z&��`   `   c�q�l�l���^���I�P�/���K�����ؾ�M��J��,������[.������,��J���M����ؾK�����P�/���I���^�l�l�`   `   A/�Ù+�.�!�
���A�X���̾�^��
[�����jۭ��ٯ��˰��ٯ�jۭ����
[���^���̾X���A�
��.�!�Ù+�`   `   ����k��F���־M�ž'A��g⭾ŵ��`]�����+����:¾�ľ�:¾+������`]��ŵ��g⭾'A��M�ž�־F��k��`   `   �ɨ��A���I��~����S������D׀���]���&˾��ھk��%��k�徍�ھ�&˾�]��׀��D�����S��~����I���A��`   `   �k���l���p��gy�o��3�����;¾�O�ھ{��6�҇����҇�6�{��O�ھ;¾���3���o���gy���p���l�`   `   P-���1���?��Y�H��O���佾+���	�'�.D1�m_=�o�A�m_=�.D1�'��	�+�澀佾O��H���Y���?���1�`   `   i������-��W����@˴�	�
��~�2���P��(i��0y���~��0y��(i���P�~�2�
��	�@˴�����W��-����`   `   ���H�F@A��h���y��R�*!��N�g�{�q	��7~������1�������7~��q	��g�{��N�*!�R�y���h��F@A��H�`   `   �&�q�'�TZ��Ř�W.پG���3L�u���ᷠ�����[��_���k��_���[����ᷠ�u����3L�G��W.پ�Ř�TZ�q�'�`   `   >r,�b3A�vv��i��s7���;��|�p����cѿ���`s*��&F�$�P��&F�`s*�����cѿp����|���;�s7�i��vv��b3A�`   `   �I���b��$���,ܾ�� ���a������˿����H�AƂ�~��1g��~��AƂ��H�����˿������a��� ��,ܾ�$����b�`   `   ��j����Yn���� ���;��X���ܥ�]*E��̏�DQ���<��,/���<��DQ���̏�]*E�ܥ���X����;��� �Yn�����`   `   �h��$�ɾc�E�T��A���.ҿ��#��s���������
P���
P���������s����#��.ҿ�A��E�T�c�$�ɾ�h��`   `   ���p�����޾�!��`h�|�����)E�秠�T����l�C�7�oA�C�7��l�T���秠�)E���|����`h��!���޾p���`   `   ����Y��w4�*V+���u�����X�p^�EV��S���g0�XHN��$Y�XHN��g0�S��EV��p^�X�������u�*V+�w4�Y��`   `   �����������)^0�͌{�?Ȱ����^g�&P���b��7�]aV���a�]aV��7��b�&P���^g���?Ȱ�͌{�)^0��������`   `   ���k���������/�jy��#��I����^�f���1��G�0��ON�w!Y��ON�G�0�1��f�����^�I���#��jy���/�����k���`   `   �Ƭ�\�����*�)�o��y��FY�$F���.����Ï7��\A�Ï7���.����$F�FY��y��)�o��*����\�`   `   ��������;����8j_��z���hտN�$�Y���d3�����<����<����d3��Y���N�$��hտ�z��8j_�����;龪��`   `   �@��,f����ھ�d���I�S�������y�O%F�����P������*��������P�����O%F�y�����S�����I��d���ھ,f��`   `   Cg���$��:�ɾ�>�1u1���n����K�οh���VH�ơ�����������ơ���VH�h��K�ο�����n�1u1��>�:�ɾ�$��`   `   �d��㵞�Ѹ�����K���I�>ۂ�~��{�ҿ9��$�)��+E�ݙO��+E�$�)�9��{�ҿ~��>ۂ���I��K����Ѹ�㵞�`   `   趐�к�������<̾�� �˜&���U�^<�����������Y������Y������������^<����U�˜&��� ��<̾����к��`   `   �K���4��;����굾5�ھ����*�7R��{��i��b�������������b����i���{�7R��*����5�ھ�굾;����4��`   `   㶑�N����m������M����޾���~!��w?�y�[��Fs��Y������Y���Fs�y�[��w?��~!����޾M��������m��N���`   `   �y��S�������F��n���3���D�־L#��dI� !��#1��;���?��;��#1� !�dI�L#��D�־3���n����F�����S���`   `   ;9�����������A�������I��q���, þC�Ծy��e���{����{��e���y��C�Ծ, þq����I�������A����������`   `   � �hs�O�ھ�̾����*4��ƨ��JK������犫�Ά��=R��-$��=R��Ά��犫�����JK��ƨ��*4�������̾O�ھhs�`   `   ��v�!��y� :�ܯȾ�ï�uJ���Ǝ�����}���/׀�)p��/׀�}��������Ǝ�uJ���ï�ܯȾ :�y�!��v�`   `   0vN�SJ��I=�H*�E0����˾x���%���k�8/P��NA�ɓ<��NA�8/P��k�%��x����˾��E0�H*��I=�SJ�`   `   ������G�{�9�a�%�A�� �Az��ҥþ�Y����i�8�;�u�!�2�u�!�8�;���i��Y��ҥþAz��� �%�A�9�a�G�{����`   `   1�������7~��q	��g�{��N�*!�R�y���h��F@A��H����H�F@A��h���y��R�*!��N�g�{�q	��7~������`   `   �k��_���[����ᷠ�u����3L�G��W.پ�Ř�TZ�q�'��&�q�'�TZ��Ř�W.پG���3L�u���ᷠ�����[��_��`   `   #�P��&F�`s*�����cѿp����|���;�s7�i��vv��b3A�>r,�b3A�vv��i��s7���;��|�p����cѿ���`s*��&F�`   `   1g��~��AƂ��H�����˿������a��� ��,ܾ�$����b��I���b��$���,ܾ�� ���a������˿����H�AƂ�~��`   `   ,/���<��DQ���̏�]*E�ܥ���X����;��� �Yn�������j����Yn���� ���;��X���ܥ�]*E��̏�DQ���<��`   `   ��
P���������s����#��.ҿ�A��E�T�c�$�ɾ�h���h��$�ɾc�E�T��A���.ҿ��#��s���������
P�`   `   oA�C�7��l�T���秠�)E���|����`h��!���޾p������p�����޾�!��`h�|�����)E�秠�T����l�C�7�`   `   �$Y�XHN��g0�S��EV��p^�X�������u�*V+�w4�Y������Y��w4�*V+���u�����X�p^�EV��S���g0�XHN�`   `   ��a�]aV��7��b�&P���^g���?Ȱ�͌{�)^0�������������������)^0�͌{�?Ȱ����^g�&P���b��7�]aV�`   `   w!Y��ON�G�0�1��f�����^�I���#��jy���/�����k������k���������/�jy��#��I����^�f���1��G�0��ON�`   `   �\A�Ï7���.����$F�FY��y��)�o��*����\��Ƭ�\�����*�)�o��y��FY�$F���.����Ï7�`   `   ���<����d3��Y���N�$��hտ�z��8j_�����;龪����������;����8j_��z���hտN�$�Y���d3�����<�`   `   *��������P�����O%F�y�����S�����I��d���ھ,f���@��,f����ھ�d���I�S�������y�O%F�����P������`   `   ������ơ���VH�h��K�ο�����n�1u1��>�:�ɾ�$��Cg���$��:�ɾ�>�1u1���n����K�οh���VH�ơ�����`   `   ݙO��+E�$�)�9��{�ҿ~��>ۂ���I��K����Ѹ�㵞��d��㵞�Ѹ�����K���I�>ۂ�~��{�ҿ9��$�)��+E�`   `   ���Y������������^<����U�˜&��� ��<̾����к��趐�к�������<̾�� �˜&���U�^<�����������Y���`   `   �������b����i���{�7R��*����5�ھ�굾;����4���K���4��;����굾5�ھ����*�7R��{��i��b������`   `   ����Y���Fs�y�[��w?��~!����޾M��������m��N���㶑�N����m������M����޾���~!��w?�y�[��Fs��Y��`   `   ��?��;��#1� !�dI�L#��D�־3���n����F�����S����y��S�������F��n���3���D�־L#��dI� !��#1��;�`   `   ��{��e���y��C�Ծ- þq����I�������A����������;9�����������A�������I��q���, þC�Ծy��e���{��`   `   -$��=R��Ά��犫�����JK��ƨ��*4�������̾O�ھhs例 �hs�O�ھ�̾����*4��ƨ��JK������犫�Ά��=R��`   `   )p��/׀�}��������Ǝ�vJ���ï�ܯȾ :�y�!��v���v�!��y� :�ܯȾ�ï�uJ���Ǝ�����}���/׀�`   `   ɓ<��NA�8/P��k�%��x����˾��E0�I*��I=�SJ�0vN�SJ��I=�I*�E0����˾x���%���k�8/P��NA�`   `   2�u�!�8�;���i��Y��ҥþAz��� �%�A�9�a�G�{����������G�{�9�a�%�A�� �Az��ҥþ�Y����i�8�;�u�!�`   `   Uo�&a"� J�KB��E���du��+�(�G�W������!��KM������¿��KM���!������G�W�+�(�du��E���KB�� J�&a"�`   `    ��L/��d�Sޟ�-�㾄9��V�T؈�yS��wο���#�
�C�#�
����wοyS��T؈��V��9�-��Sޟ��d��L/�`   `   �84�q�I��^���������sE���������$�@>���=��^�)[j��^���=�@>��$῰������sE���������^��p�I�`   `   ��R��m��&��n��s(���l�Hw���ڿũ�#�`�ث��$���q̸�$���ث��#�`�ũ��ڿHw����l�s(�n���&���m�`   `   ��t�Xى�.�����zE�k����Ծ�k-��T]�o���tj�����*�����tj��o����T]�k-��Ծ�k���zE���.���Xى�`   `   �k���Ɯ�)�Ҿ�~��^�dӛ�uC⿁%6��r��#V��|��Y)���2��Y)�|�#V���r���%6�uC�dӛ��^��~�)�Ҿ�Ɯ�`   `   �t���a������(��ds�x���?��8S]�����o�*-0��N��X��N�*-0��o����7S]�?��x����ds���(��辏a��`   `   2��c���o��Ea3����
ƶ�9��z�y��	��5F��<g�̄s��<g��5F�	�y���z�9�
ƶ����Ea3��o��c��`   `   >�������/ �ra8����F��@;�\���h��#\��N��\p��m}��\p��N�#\��h��\��@;�F�����ra8�/ �����`   `   ����5ľ�� �pt7�U���#��n���tz�ޢ�����CF�v@g���s�v@g��CF���ޢ���tz�n���#��U��pt7��� ��5ľ`   `   V"��Ł���$���0�i-z�4H��k��8^�P6��\���=0�}N�t�X�}N��=0�\��P6��8^�k��4H��i-z��0��$��Ł��`   `   )쩾�u��vF�t%��h��Ο��J忩97�&Γ�����W�>O)�~�2�>O)�W�����&Γ��97��J忬Ο��h�t%�vF��u��`   `   Q����B���ܾC���Q�������¿�w��^�-ڢ��i���x���o��x���i��-ڢ��^��w���¿�����Q�C���ܾ�B��`   `   T����k���Tɾ���[�7�ix������nݿ=g�?�`����� s��Y�� s������?�`�=g��nݿ����ix�[�7�����Tɾ�k��`   `   �\��ݰ���ȵ����j����Q�m����L���[⿯>��u=�"V]��wi�"V]��u=��>��[⿕L��m�����Q�j����龐ȵ�ݰ��`   `   ���x��ƹ��c�˾�m�)i,���^�gF�����W�Ϳ�9��U�	���U�	��9��W�Ϳ���gF����^�)i,��m�c�˾ƹ��x��`   `   ����׉� ���j�����ܾ�����0���[�򛃿��������阹��۾�阹���������򛃿��[���0������ܾj��� ����׉�`   `   �.��]ދ����&���k�����㾔�
�2�(�1aH�QUf�:�~�'����s��'���:�~�QUf�1aH�2�(���
����k���&������]ދ�`   `   �r������	�����a����qݾ@� �7��B�(���9��E��I��E���9�B�(�7��@� ��qݾa�����	������r���`   `   G���紾e�䮾���x���)󺾵9ʾ��ݾ(^��R��
��j��
��R�(^��ݾ�9ʾ)�x�������䮾e�紾`   `   ���p澯�ܾL�Ͼ���C���6­��4���w�����ǯ��]龾T���]龾ǯ������w���4��6­�C������L�Ͼ��ܾp�`   `   M��;����p���B쾖.Ͼ#յ���lz���[���O��󹆾�Z��󹆾�O���[��lz����#յ��.Ͼ�B�p������;�`   `   3oV�@�Q�=�D���0��!� ��Ӿ r��Lˏ� u��dY�<J�n/E�<J��dY� u�Lˏ� r���Ӿ!� ����0�=�D�@�Q�`   `   \���%d��4h��Ҫk��PJ�Ua&�����I̾}蜾��s�-PD��)�a5 ��)�-PD���s�}蜾�I̾���Ua&��PJ�Ҫk�4h��%d��`   `   ��¿��KM���!������G�W�+�(�du��E���KB�� J�&a"�Uo�&a"� J�KB��E���du��+�(�G�W������!��KM����`   `   C�#�
����wοyS��T؈��V��9�-��Sޟ��d��L/� ��L/��d�Sޟ�-�㾃9��V�T؈�yS��wο���#�
�`   `   )[j��^���=�@>��$῰������sE���������^��q�I��84�q�I��^���������sE���������$�@>���=��^�`   `   q̸�$���ث��#�`�ũ��ڿHw����l�s(�n���&���m���R��m��&��n��s(���l�Hw���ڿũ�#�`�ث��$���`   `   *�����tj��o����T]�k-��Ծ�k���zE���.���Xى���t�Xى�.�����zE�k����Ծ�k-��T]�o���tj�����`   `   ��2��Y)�|�#V���r���%6�uC�dӛ��^��~�)�Ҿ�Ɯ��k���Ɯ�)�Ҿ�~��^�dӛ�uC⿁%6��r��#V��|��Y)�`   `   �X��N�*-0��o����7S]�?��x����ds���(��辏a���t���a������(��ds�x���?��7S]�����o�*-0��N�`   `   ̄s��<g��5F�	�y���z�9�
ƶ����Ea3��o��c��2��c���o��Ea3����
ƶ�9��z�y��	��5F��<g�`   `   �m}��\p��N�#\��h��\��@;�F�����ra8�/ �����>�������/ �ra8����F��@;�\���h��#\��N��\p�`   `   ��s�v@g��CF���ޢ���tz�n���#��U��pt7��� ��5ľ����5ľ�� �pt7�U���#��n���tz�ޢ�����CF�v@g�`   `   t�X�}N��=0�\��P6��8^�k��4H��i-z��0��$��Ł��V"��Ł���$���0�i-z�4H��k��8^�P6��\���=0�}N�`   `   ~�2�>O)�W�����&Γ��97��J忬Ο��h�t%�vF��u��)쩾�u��vF�t%��h��Ο��J忩97�&Γ�����W�>O)�`   `   �o��x���i��-ڢ��^��w���¿�����Q�C���ܾ�B��Q����B���ܾC���Q�������¿�w��^�-ڢ��i���x��`   `   Y�� s������?�`�=g��nݿ����ix�[�7�����Tɾ�k��T����k���Tɾ���[�7�ix������nݿ=g�?�`����� s��`   `   �wi�"V]��u=��>��[⿕L��m�����Q�j����龐ȵ�ݰ���\��ݰ���ȵ����j����Q�m����L���[⿯>��u=�"V]�`   `   ��U�	��9��W�Ϳ���gF����^�)i,��m�c�˾ƹ��y�����y��ƹ��c�˾�m�)i,���^�gF�����W�Ϳ�9��U�	�`   `   �۾�阹���������򛃿��[���0������ܾk��� ����׉�����׉� ���k�����ܾ�����0���[�򛃿��������阹�`   `   �s��'���:�~�QUf�1aH�2�(���
����k���&������]ދ��.��]ދ����&���k�����㾔�
�2�(�1aH�QUf�:�~�'���`   `   �I��E���9�B�(�7��@� ��qݾa�����	������r����r������	�����a����qݾ@� �7��B�(���9��E�`   `   �j��
��R�(^��ݾ�9ʾ)�x�������䮾e�紾G���紾e�䮾���x���)󺾵9ʾ��ݾ(^��R��
�`   `   T���]龾ǯ������w���4��6­�C������L�Ͼ��ܾp����p澯�ܾL�Ͼ���C���6­��4���w�����ǯ��]龾`   `   �Z��󹆾�O���[��lz����#յ��.Ͼ�B�p������;�M��;����p���B쾖.Ͼ#յ���lz���[���O��󹆾`   `   n/E�<J��dY� u�Lˏ� r���Ӿ!� ����0�=�D�@�Q�3oV�@�Q�=�D���0��!� ��Ӿ r��Lˏ� u��dY�<J�`   `   a5 ��)�-PD���s�}蜾�I̾���Ua&��PJ�Ҫk�4h��%d��\���%d��4h��Ҫk��PJ�Ua&�����I̾}蜾��s�-PD��)�`   `   �8�9;#��K��������g���}�)���X��M��s��h��
e��Ŀ
e��h��s���M����X�}�)�g�����������K�9;#�`   `   ����80�ZJe�����$��a �?5W�N���<f��!п�N��ff�1��ff��N��!п<f��N���?5W�a �$�侢���ZJe��80�`   `   �(5�`K�_��Y�����)&F�T̄������*���j@�~)a�|�m�~)a�j@����*㿇���T̄�)&F���Y���_��`K�`   `   P�S�6@n�����/��g)��m��p����ܿ#��K�c��Ε�P=���|��P=���Ε�K�c�#����ܿ�p���m��g)�/�����6@n�`   `   �/v�F���Q������D#F�[v��@�����vi`�{��W���^&��y�^&�W���{��vi`����@��[v��D#F����Q���F���`   `   �������O
Ծ�Z�0�_���T�=�8�����/������+��5��+���/�������<�8��T��0�_��Z�O
Ծ����`   `   I)��5�����{�)��t�F���7!��g`������`��2�.�P���[�.�P��2��`������g`�7!�F����t�{�)����5��`   `   �妾
캾8���+[4�7T���
�����g�}�3����2���H��]j���v��]j���H��2�3���g�}�����
��7T��+[4�8���
캾`   `   XV����¾���Z9�9I���������8�������� ���P�Y�s�|���Y�s���P��� ������8��������9I���Z9�����¾`   `   !���ľr�&c8� ���e��L@���}����nB�y�H�9aj�F�v�9aj�y�H�nB������}�L@��e�� ��&c8�r��ľ`   `   �|��� ¾����1��s{��b���)��%a�8ݸ��x�'�2���P���[���P�'�2��x�8ݸ��%a��)��b���s{��1����� ¾`   `   �	��V�����)&�,�i������U�D�9�������@�]�+���4�]�+�@�������D�9��U翔���,�i��)&����V���`   `   �С��<���Tݾ_��R�{����ÿ��'a�Z8��ɏ���6a��ɏ��Z8��'a�����ÿ{���R�_��Tݾ�<��`   `   ))�����eɾ��R8�`�y�����S߿bL ���c�P������7����P�����c�bL ��S߿���`�y�R8����eɾ��`   `   ����)��䎵�R0�_���R��?���f��+^�1����?��j`��l��j`���?�1��+^��f���?����R�_�R0�䎵�)��`   `   �B��HM���F��a�˾G��%-�g�_�������dzϿ̢��y8��c�y8�̢��dzϿ������g�_�%-�G��a�˾�F��HM��`   `   =3�����/ ���d��BZݾ��z�1�/�\��O���~��G�����G����G����~���O��/�\�z�1���BZݾ�d��/ �����`   `   �T����[����z��f������R�])��tI�c�g����R��:���R����c�g��tI�])�R����f����z��[�����`   `   \O��� ���"��$֡�5���¾�M޾`'�ǉ�q�)�O�:��2F��-J��2F�O�:�q�)�ǉ�`'��M޾�¾5��$֡��"��� ��`   `   Tߵ������ձ�w��P��]������˾�߾«��R���
�46���
�R�«���߾�˾���]���P��w󮾙ձ�����`   `   �4꾮��3\ݾоW¾��g���﫾*J�����e����򿾈�����e������*J���﫾g����W¾о3\ݾ���`   `   ���D��c�bV��)� о�����͢�,��������xo��r��xo��������,���͢������ о�)�bV�c�D��`   `   �lW���R��E���1���Q$�֪Ծ�D���|���Pv��Z�[K��7F�[K��Z��Pv��|���D��֪ԾQ$�����1��E���R�`   `   �M�����}����l�`K�oC'�����V;#���a�t��RE�|�)��!�|�)��RE�a�t�#����V;���oC'�`K���l�}�����`   `   Ŀ
e��h��s���M����X�}�)�g�����������K�9;#��8�9;#��K��������g���}�)���X��M��s��h��
e��`   `   1��ff��N��!п<f��N���?5W�a �$�侢���ZJe��80�����80�ZJe�����$��a �?5W�N���<f��!п�N��ff�`   `   {�m�~)a�j@����*㿇���T̄�)&F���Y���_��`K��(5�`K�_��Y�����)&F�T̄������*���j@�~)a�`   `   �|��P=���Ε�K�c�#����ܿ�p���m��g)�/�����6@n�P�S�6@n�����/��g)��m��p����ܿ#��K�c��Ε�P=��`   `   �y�^&�W���{��vi`����@��[v��D#F����Q���F����/v�F���Q������D#F�[v��@�����vi`�{��W���^&�`   `   �5��+���/�������<�8��T��0�_��Z�O
Ծ�����������O
Ծ�Z�0�_���T�<�8�����/������+�`   `   ��[�.�P��2��`������g`�7!�F����t�{�)����5��I)��5�����{�)��t�F���7!��g`������`��2�.�P�`   `   ��v��]j���H��2�3���g�}�����
��7T��+[4�8���
캾�妾
캾8���+[4�7T���
�����g�}�3����2���H��]j�`   `   |���Y�s���P��� ������8��������9I���Z9�����¾XV����¾���Z9�9I���������8�������� ���P�Y�s�`   `   F�v�9aj�y�H�nB������}�L@��e�� ��&c8�r��ľ!���ľr�&c8� ���e��L@���}����nB�y�H�9aj�`   `   ��[���P�'�2��x�8ݸ��%a��)��b���s{��1����� ¾�|��� ¾����1��s{��b���)��%a�8ݸ��x�'�2���P�`   `   ��4�]�+�@�������D�9��U翔���,�i��)&����V����	��V�����)&�,�i������U�D�9�������@�]�+�`   `   6a��ɏ��Z8��'a�����ÿ{���R�_��Tݾ�<���С��<���Tݾ_��R�{����ÿ��'a�Z8��ɏ���`   `   �7����P�����c�bL ��S߿���`�y�R8����eɾ��))�����eɾ��R8�`�y�����S߿bL ���c�P�����`   `   �l��j`���?�1��+^��f���?����R�_�R0�厵�)������)��厵�R0�_���R��?���f��+^�1����?��j`�`   `   �c�y8�̢��dzϿ������g�_�%-�G��b�˾�F��HM���B��HM���F��b�˾G��%-�g�_�������dzϿ̢��y8�`   `   G����G����~���O��/�\�z�1���BZݾ�d��/ �����>3�����/ ���d��BZݾ��z�1�/�\��O���~��G�����`   `   :���R����c�g��tI�])�R����f����z��[�������T�����[����z��f������R�])��tI�c�g����R��`   `   �-J��2F�O�:�q�)�ǉ�`'��M޾�¾5��$֡��"��� ��\O��� ���"��$֡�5���¾�M޾`'�ǉ�q�)�O�:��2F�`   `   46���
�R�«���߾�˾���]���P��w󮾙ձ�����Tߵ������ձ�w��P��]������˾�߾«��R���
�`   `   ������e������*J���﫾g����W¾о3\ݾ����4꾮��3\ݾоW¾��g���﫾*J�����e�����`   `   r��xo��������,���͢������ о�)�cV�d�D�����D��d�cV��)� о�����͢�,��������xo��`   `   �7F�[K��Z��Pv��|���D��֪ԾQ$�����1��E���R��lW���R��E���1���Q$�֪Ծ�D���|���Pv��Z�[K�`   `   �!�|�)��RE�a�t�#����V;���oC'�`K���l�}������M�����}����l�`K�oC'�����V;#���a�t��RE�|�)�`   `   �)����KD�q���M��C���y�#�9|Q�?��4y���|���9���Q���9���|��4y��?��9|Q�y�#�C����M��q���KD���`   `   ����O*��]� =��Q�ܾ�]�q�O�`Ȅ�������ſ���D�u��D���鿞�ſ����`Ȅ�q�O��]�Q�ܾ =���]��O*�`   `   �(/��?D�����V��>}��?�I"������0�ֿ�D��0��2N�HZY��2N��0��D�0�ֿ����I"���?�>}�V�������?D�`   `   �L�nf�p����߾�D#�{�e��G��øпo���GP��x��BR��5���BR���x���GP�o��øп�G��{�e��D#��߾p���nf�`   `   gn�����C��S��
?������g�����@EM��*�������7������7�������*��@EM�����g������
?�S���C�����`   `   �Շ�띘�G�̾D��DX��ږ�O�׿)�)�	-���s��_����){%����_��s��	-��)�)�O�׿�ږ�DX�D��G�̾띘�`   `   ����������ж#�^5l�򤥿3���CM�Pק�R��()#�@?��tI�@?�()#�R��Pק��CM�3��򤥿^5l�ж#��⾍���`   `   �|��U��� ��.�F�y����b���qg�:�������7���V�b���V��7����:����qg�b�����F�y��.� ��U���`   `   OP��Ͱ��jv��s#3����mU���A�Y>q�H���ށ��??�d,_��j�d,_��??�ށ�H���Y>q��A�lU�����s#3�jv��Ͱ��`   `   "譾I��������w2�}O}������+�u�g�B���=��!�7�f�V�}	b�f�V�!�7�=��B���u�g��+�����}O}��w2�����I���`   `   �}�����HE���g,��Ts��w���m��0/N��@�������E#��??�ceI��??��E#������@��0/N��m���w���Ts��g,�HE�����`   `   X����j����ս!�֞b�����1�ڿ��*�ť��}����)�ּ��Y%�ּ��)�}���ť����*�1�ڿ����֞b�ս!��꾬j��`   `   �E��Ұ��?۾�����L�$Њ�iM���3�\0N�Fj��F��������R������F���Fj��\0N��3�iM��$Њ���L�����?۾Ұ�`   `   A�������nɾ���3���q�+���Ȝӿ^���P�W������4������W���P�^��Ȝӿ+�����q���3���nɾ���`   `   ᭓��[��r����o�F��'�L�@ф�o{����׿�D�!p0��FM��HX��FM�!p0��D���׿o{��@ф�'�L�F���o�r����[��`   `   �n��?Ǔ�㹧�;�˾��v�(���X��Q���i���<ſ��翂��U9������翸<ſ�i���Q����X�v�(���;�˾㹧�?Ǔ�`   `   �͊�����\���ാ=E۾A��!o,��rU����⓿d���ϝ��En��ϝ��d����⓿���rU�!o,�A��=E۾�ാ�\�����`   `   �s���������>i���׽�)y�@����#��B�i�_�DKw�P����E��P���DKw�i�_��B���#�@��(yྷ׽�>i���������`   `   �]���D���J��A��������ؾ���D���#��$4��?���B��?��$4��#�D�������ؾ���A����J���D��]��`   `   �緾z}���鲾��������Y���o��/xž�ؾdW쾚���i����i������dW쾛ؾ/xž�o���Y����������鲾z}��`   `   t�����F۾N�;���~���Ea���P������#��|Z���L���,���L��|Z���#������P��Ea��~������N�;�F۾���`   `   �v�sn�����O�}�羳�ʾձ�H��L���l���'���`₾R~��`₾'���l���L���H��ձ���ʾ}���O����sn�`   `   �/Q���L���?�o,�N7�����Mξk�������n��aS��YD��?��YD��aS���n����k���Mξ���N7�o,���?���L�`   `   �������e���+e�
�D��!��3 ��ƾ����m�^�>�UF$�I��UF$�^�>��m�����ƾ�3 ��!�
�D��+e�e������`   `   �Q���9���|��4y��?��9|Q�y�#�C����M��q���KD����)����KD�q���M��C���y�#�9|Q�?��4y���|���9��`   `   u��D���鿞�ſ����`Ȅ�q�O��]�Q�ܾ =���]��O*�����O*��]� =��Q�ܾ�]�q�O�`Ȅ�������ſ���D�`   `   HZY��2N��0��D�/�ֿ����I"���?�>}�V�������?D��(/��?D�����V��>}��?�I"������/�ֿ�D��0��2N�`   `   5���AR���x���GP�o��øп�G��{�e��D#��߾p���nf��L�nf�p����߾�D#�{�e��G��øпo���GP��x��AR��`   `   ����7�������*��@EM�����g������
?�S���C�����gn�����C��S��
?������g�����@EM��*�������7��`   `   ){%����_��s��	-��)�)�O�׿�ږ�DX�D��G�̾띘��Շ�띘�G�̾D��DX��ږ�O�׿)�)�	-���s��_����`   `   �tI�@?�()#�R��Pק��CM�3��򤥿^5l�ж#��⾍�������������ж#�^5l�򤥿3���CM�Pק�R��()#�@?�`   `   b���V��7����:����qg�b�����F�y��.� ��U����|��U��� ��.�F�y����b���qg�:�������7���V�`   `   �j�d,_��??�ށ�H���Y>q��A�mU�����s#3�jv��Ͱ��OP��Ͱ��jv��s#3����mU���A�Y>q�H���ށ��??�d,_�`   `   }	b�f�V�!�7�=��B���u�g��+�����}O}��w2�����I���"譾I��������w2�}O}������+�u�g�B���=��!�7�f�V�`   `   ceI��??��E#������@��0/N��m���w���Ts��g,�HE������}�����HE���g,��Ts��w���m��0/N��@�������E#��??�`   `   �Y%�ּ��)�}���ť����*�1�ڿ����֞b�ս!��꾬j��Y����j����ս!�֞b�����1�ڿ��*�ť��}����)�ּ�`   `   �R������F���Fj��\0N��3�iM��$Њ���L�����?۾Ұ��E��Ұ��?۾�����L�$Њ�iM���3�\0N�Fj��F�������`   `   4������W���P�^��Ȝӿ+�����q���3���nɾ���A�������nɾ���3���q�+���Ȝӿ^���P�W������`   `   �HX��FM�!p0��D���׿o{��@ф�'�L�F���o�r����[��⭓��[��r����o�F��'�L�@ф�o{����׿�D�!p0��FM�`   `   U9������翸<ſ�i���Q����X�v�(���;�˾㹧�?Ǔ��n��?Ǔ�㹧�;�˾��v�(���X��Q���i���<ſ��翂��`   `   En��ϝ��d����⓿���rU�!o,�A��=E۾�ാ�\������͊�����\���ാ=E۾A��!o,��rU����⓿d���ϝ��`   `   �E��Q���DKw�i�_��B���#�@��)yྷ׽�>i����������s���������>i���׽�)y�@����#��B�i�_�DKw�Q���`   `   ��B��?��$4��#�E�������ؾ���A����J���D��]���]���D���J��A��������ؾ���D���#��$4��?�`   `   ��i������dW쾛ؾ/xž�o���Y����������鲾z}���緾z}���鲾��������Y���o��/xž�ؾdW쾚���i��`   `   �,���L��|Z���#������P��Ea��~������N�;�F۾���t�����F۾N�;���~���Ea���P������#��|Z���L��`   `   R~��`₾'���l���L���H��ձ���ʾ}���O����sn��v�sn�����O�}�羳�ʾձ�H��L���l���'���`₾`   `   �?��YD��aS���n����k���Mξ���N7�o,���?���L��/Q���L���?�o,�N7�����Mξk�������n��aS��YD�`   `   I��UF$�^�>��m�����ƾ�3 ��!�
�D��+e�e�������������e���+e�
�D��!��3 ��ƾ����m�^�>�UF$�`   `   T��!|�x6�ryt�뇧�� �4��9B�tim�����ug��:��U��:��ug������tim�9B�4��� �뇧�ryt�x6�!|�`   `   ����,���M�����x̾���+@�v������Z���oϿ/b���/b��oϿ�Z������v�+@�����x̾�����M��,�`   `   $�"�m6�Air��Z��jg���0�sEm��;���H��v��g��,�I�4��,�g�v���H���;��sEm��0�jg���Z��Air�m6�`   `   ��>���V�y���t0Ͼ����eT�GD��m��M���AY-��(`�d��~q��d���(`�AY-�M���m��GD���eT����t0Ͼy�����V�`   `   Դ^��"z�s~��o[�}0�1.w�� ��$����*�N�u����U޿�R���U޿����N�u���*�$�迋 ��1.w�}0�o[�s~���"z�`   `   ̪~�����d���T�	���G�uC��l������`_�U���@��Fg �H��Fg ��@��U��`_����l���uC����G�T�	�d�������`   `   G�����a�Ҿ��<�Z�9���&ٿ��*����l��5���p�#&��p�5���l������*��&ٿ9��<�Z���a�Ҿ����`   `   N��G����}�!�y�g�R2��Rz�HR?��?������~"��q1�;��q1�~"������?��HR?�Rz�R2��y�g�}�!��G���`   `   ������J�뾋�&��am��礿���hG����z���mp�z�8�npB�z�8�mp�z������hG����礿�am���&�J�����`   `   M���?���5����&���k��ʢ�E���?�E���E���E�{1�x ;�{1�E�E���E����?�E�쿛ʢ���k���&�5��?���`   `   .b��6	���0�~F"�$c�<c��Q�ۿ' ,�Z���c������op��&�op����c���Z���& ,�Q�ۿ<c��$c�~F"��0�6	��`   `   	���#Y��"�����5hT���;Ŀx���`����hu���M �����M �hu������`�x���;Ŀ�5hT����"��#Y��`   `   �����S���ھ�N�p A�����R�����,�?av�f��*|��Jm��*|��f��?av�,����R������p A��N��ھ�S��`   `   ����%ͯ��%;�\���*��c��>��؟��Ω����-���_��r���Ҋ��r����_���-�Ω��؟���>���c���*��\��%;%ͯ�`   `   |���?�������`�(��A�A"x��f�������������*�pc3���*�����������f��A"x��A�(��`����?���`   `   U��,��*P����Ͼ���fI �=K�x�{���������oͿ>�⿯��>�⿓oͿ�������x�{�=K�fI ������Ͼ*P��,��`   `   ]������~���Oƻ��	ھ���M"���F��lm�҈��?��x�����x���?��҈��lm���F��M"����	ھOƻ�~������`   `   �A��XF��+'�����
s7ھ�� �7�͡4�� O�e� ts�Q�x� ts�e�� O�͡4�7��� �s7ھ
���+'��XF��`   `   :�������Ѩ�����������wdϾ�������N�&���0�4���0�N�&��������wdϾ�����������Ѩ�����`   `   �F���1�������������u����
���Aʾ{�۾����f��$����f�����{�۾Aʾ
������u�������������1��`   `   �d�̕��
ھ�%˾'��}�������u��3����u�����SΫ�hm��SΫ�����u��3����u�����}���'���%˾�
ھ̕�`   `   (�����h�	�/K����ݾl���#ܨ��~����u^��v�}8s��Rr�}8s��v�u^����~��#ܨ�l�����ݾ/K��h�	����`   `   pTE��A���4�M"�Z���k���E����7���^���D�"�6�^�1�"�6���D��^��7��E���k�����Z�M"���4��A�`   `   bf������n���U��7��o�M��#=���d����\�/�1�a��H}�a��/�1���\��d��#=��M�o��7���U���n���`   `   U��:��ug������tim�9B�4��� �뇧�ryt�x6�!|�T��!|�x6�ryt�뇧�� �4��9B�tim�����ug��:��`   `   ��/b��oϿ�Z������v�+@�����x̾�����M��,�����,���M�����x̾���+@�v������Z���oϿ/b�`   `   I�4��,�g�v���H���;��sEm��0�jg���Z��Air�m6�$�"�m6�Air��Z��jg���0�sEm��;���H��v��g��,�`   `   ~q��d���(`�AY-�M���m��GD���eT����t0Ͼy�����V���>���V�y���t0Ͼ����eT�GD��m��M���AY-��(`�d��`   `   R���U޿����N�u���*�$�迋 ��1.w�}0�o[�s~���"z�Դ^��"z�s~��o[�}0�1.w�� ��$����*�N�u����U޿�`   `   H��Fg ��@��U��`_����l���uC����G�T�	�d�������̪~�����d���T�	���G�uC��l������`_�U���@��Fg �`   `   #&��p�5���l������*��&ٿ9��<�Z���a�Ҿ����G�����a�Ҿ��<�Z�9���&ٿ��*����l��5���p�`   `   ;��q1�~"������?��HR?�Rz�R2��y�g�}�!��H���N��H����}�!�y�g�R2��Rz�HR?��?������~"��q1�`   `   npB�z�8�mp�z������hG����礿�am���&�J�����������J�뾋�&��am��礿���hG����z���mp�z�8�`   `   x ;�{1�E�E���E����?�E�쿛ʢ���k���&�5��?���M���?���5����&���k��ʢ�E���?�E���E���E�{1�`   `   �&�op����c���Z���& ,�Q�ۿ<c��$c�~F"��0�6	��.b��6	���0�~F"�$c�<c��Q�ۿ& ,�Z���c������op�`   `   ����M �hu������`�x���;Ŀ�5hT����"��#Y��
���#Y��"�����5hT���;Ŀx���`����hu���M �`   `   Jm��*|��f��?av�,����R������p A��N��ھ�S�������S���ھ�N�p A�����R�����,�?av�f��*|��`   `   �Ҋ��r����_���-�Ω��؟���>���c���*��\��%;%ͯ�����%ͯ��%;�\���*��c��>��؟��Ω����-���_��r��`   `   pc3���*�����������f��A"x��A�(��`����?���|���?�������`�(��A�A"x��f�������������*�`   `   ���>�⿓oͿ�������x�{�=K�fI ������Ͼ*P��,��U��,��*P����Ͼ���fI �=K�x�{���������oͿ>��`   `   ���x���?��҈��lm���F��M"����	ھOƻ�������]���������Oƻ��	ھ���M"���F��lm�҈��?��x��`   `   Q�x� ts�e�� O�͡4�7��� �s7ھ
���+'��XF���A��XF��+'�����
s7ھ�� �7�͡4�� O�e� ts�`   `   4���0�N�&��������wdϾ�����������Ѩ�����:�������Ѩ�����������wdϾ�������N�&���0�`   `   $����f�����|�۾Aʾ
������u�������������1���F���1�������������u����
���Aʾ{�۾����f��`   `   hm��SΫ�����u��3����u�����}���'���%˾�
ھ̕依d�̕��
ھ�%˾'��}�������u��3����u�����SΫ�`   `   �Rr�}8s��v�u^����~��#ܨ�l�����ݾ/K��h�	����(�����h�	�/K����ݾl���#ܨ��~����u^��v�}8s�`   `   ^�1�"�6���D��^��7��E���k�����Z�M"���4��A�pTE��A���4�M"�Z���k���E����7���^���D�"�6�`   `   H}�a��/�1���\��d��#=��M�o��7���U���n���bf������n���U��7��o�M��#=���d����\�/�1�a��`   `   ���(��k#���Z����K�˾�9��3-��KT��Cx�EȊ�ƌ�� ��ƌ��EȊ��Cx��KT��3-��9�K�˾�����Z�k#�(��`   `   ���3���7�����q���T6��.`*��Z�߅���&���p���8ǿ�p��&����߅��Z�.`*�T6��q���������7�3�`   `   ���y#�-iX��L��g�ݾ�%���R�Ć�UP��ǚɿ���	.����	.����ƚɿUP��Ć���R��%�g�ݾ�L��-iX�y#�`   `   �}+�#i@�eI���'���^�<�;|��n��K�п ����(��D�}}N��D���(� ��K�п�n��;|�<��^��'��eI��#i@�`   `   �?I�ma������X׾�#��B[������+¿��_@7���m��D���M���D����m�_@7����+¿�����B[��#��X׾����ma�`   `   ��g��r��n4�������1�=w��O��e�Q�'�w�p�����i����v��i�������w�p�Q�'�e��O��=w��1�����n4���r��`   `   j���%���B��4�CYB�����<ɷ�J����J�H����X����O:�����X��H�����J�J��<ɷ�����CYB�4��B��%��`   `   U㏾F螾��;g��{YN��^��^tĿ����9d�Z����x��0��
�0���x��Z����9d����^tĿ�^��{YN�g����;F螾`   `   8d��;O���پ_d��DT�1���;�ɿa��^�m��߮�����9�^���9�����߮�^�m�a��;�ɿ1����DT�_d��پ;O��`   `   �K���u�� �߾��-�S�*]��K�ſ�=���d�)����������
��������)����d��=�K�ſ*]��-�S��� �߾�u��`   `   ����Q���$㾹4���M��Ċ�����,���K�M��ٰ����������ٰ��M����K�,������Ċ���M��4�$�Q���`   `   嫵�����+"�"U��WB�Ԝ���~��<�7I)���q������g������g��������q�7I)�<鿚~��Ԝ���WB�"U�+"㾢���`   `   Fv���ž���VT
�ZK3��uk����w�ſ�,�Q�7��m�7ߋ�r���7ߋ��m�Q�7��,�w�ſ����uk�ZK3�VT
�����ž`   `   �¾�VȾX�ܾ<	�v"��P�����sJ��+�ҿ���h(�}C��/M�}C��h(���+�ҿsJ�������P�v"�<	�X�ܾ�VȾ`   `   ƾz�ɾR׾�Z�X��M3�Ea��Ǌ����a�ɿ�-�'��ԅ
�'���-�a�ɿ����Ǌ�Ea��M3�X��Z�R׾z�ɾ`   `   c�Ǿ��ɾ��оb��X��������9���b�����5������#���ÿ�#������5�������b���9����X���b�ྜ�о��ɾ`   `   �_ȾmȾ��ɾ۔о�������;�ԭ3�NOT�k�s��ǆ�����5��������ǆ�k�s�NOT�ԭ3��;�������۔о��ɾmȾ`   `   z�ȾmǾ�ľz�þ��Ⱦ	l׾���ٕ�~�!��=8��JK���W��n\���W��JK��=8�~�!�ٕ����	l׾��Ⱦz�þ�ľmǾ`   `   't̾e�ɾj�þ{���e��	ͺ��ž�پj��1@����0�;�0����0@�j���پ�ž	ͺ��e��{��j�þe�ɾ`   `   �9ؾ�Ծ-B˾8���������vĨ�+����㷾C'ž�Ҿ,�۾[�޾,�۾�ҾC'ž�㷾+���vĨ�������8���-B˾�Ծ`   `    ^�1�����n�ξ�˺��ۨ��s��K���R7��'����
��#��E^��#���
��'���R7��K����s���ۨ��˺�n�ξ���1��`   `   !�O��f��|�ZԾ𐷾uW��6s���x��$g���]��cY��@X��cY���]��$g��x�6s��uW��𐷾�ZԾ�|�f�O�`   `   xk7�|O3���'��:�ˢ��پ.)���2����n��ZI���0�i##�Z��i##���0��ZI���n��2��.)���پˢ��:���'�|O3�`   `   ��l�+�g��bX��LA��9%����ҍ׾�H���z����F����/��� ��/�����F��z���H��ҍ׾����9%��LA��bX�+�g�`   `    ��ƌ��EȊ��Cx��KT��3-��9�K�˾�����Z�k#�(�����(��k#���Z����K�˾�9��3-��KT��Cx�EȊ�ƌ��`   `   �8ǿ�p��&����߅��Z�.`*�T6��q���������7�4����4���7�����q���T6��.`*��Z�߅���&���p��`   `   ���	.����ƚɿUP��Ć���R��%�g�ݾ�L��-iX�y#����y#�-iX��L��g�ݾ�%���R�Ć�UP��ƚɿ���	.�`   `   }}N��D���(� ��K�п�n��;|�<��^��'��eI��#i@��}+�#i@�eI���'���^�<�;|��n��K�п ����(��D�`   `   �M���D����m�_@7����+¿�����B[��#��X׾����ma��?I�ma������X׾�#��B[������+¿��_@7���m��D��`   `   �v��i�������w�p�Q�'�e��O��=w��1�����n4���r����g��r��n4�������1�=w��O��e�Q�'�w�p�����i���`   `   O:�����X��H�����J�J��<ɷ�����CYB�4��B��%��j���%���B��4�CYB�����<ɷ�J����J�H����X����`   `   
�0���x��Z����9d����^tĿ�^��{YN�g����;F螾U㏾F螾��;g��{YN��^��^tĿ����9d�Z����x��0��`   `   ^���9�����߮�^�m�a��;�ɿ1����DT�_d��پ;O��8d��;O���پ_d��DT�1���;�ɿa��^�m��߮�����9�`   `   �
��������)����d��=�K�ſ*]��-�S��� �߾�u���K���u�� �߾��-�S�*]��K�ſ�=���d�)���������`   `   �����ٰ��M����K�,������Ċ���M��4�$�Q�������Q���$㾹4���M��Ċ�����,���K�M��ٰ�����`   `   ����g��������q�7I)�<鿚~��Ԝ���WB�"U�+"㾢���嫵�����+"�"U��WB�Ԝ���~��<�7I)���q������g��`   `   r���8ߋ��m�Q�7��,�w�ſ����uk�ZK3�VT
�����žFv���ž���VT
�ZK3��uk����w�ſ�,�Q�7��m�8ߋ�`   `   �/M�}C��h(���+�ҿsJ�������P�v"�<	�X�ܾ�VȾ�¾�VȾX�ܾ<	�v"��P�����sJ��+�ҿ���h(�}C�`   `   ԅ
�'���-�a�ɿ����Ǌ�Ea��M3�X��Z�R׾z�ɾƾz�ɾR׾�Z�X��M3�Ea��Ǌ����a�ɿ�-�'��`   `   �ÿ�#������5�������b���9����X���b�ྜ�о��ɾc�Ǿ��ɾ��оb��X��������9���b�����5������#��`   `   5��������ǆ�k�s�NOT�ԭ3��;�������۔о��ɾmȾ�_ȾmȾ��ɾ۔о�������;�ԭ3�NOT�k�s��ǆ�����`   `   �n\���W��JK��=8�~�!�ٕ����	l׾��Ⱦz�þ�ľmǾ{�ȾmǾ�ľz�þ��Ⱦ	l׾���ٕ�~�!��=8��JK���W�`   `   ;�0����1@�j���پ�ž	ͺ��e��	{��j�þe�ɾ't̾e�ɾj�þ{���e��	ͺ��ž�پj��1@����0�`   `   [�޾,�۾�ҾD'ž�㷾+���vĨ�������8���-B˾�Ծ�9ؾ�Ծ-B˾8���������vĨ�+����㷾C'ž�Ҿ,�۾`   `   E^��#���
��'���R7��K����s���ۨ��˺�n�ξ���1�� ^�1�����n�ξ�˺��ۨ��s��K���R7��'����
��#��`   `   �@X��cY���]��$g��x�6s��uW��𐷾�ZԾ�|�f�O�!�O��f��|�ZԾ𐷾uW��6s���x��$g���]��cY�`   `   Z��i##���0��ZI���n��2��.)���پˢ��:���'�|O3�xk7�|O3���'��:�ˢ��پ.)���2����n��ZI���0�i##�`   `   �� ��/�����F��z���H��ҍ׾����9%��LA��bX�,�g���l�,�g��bX��LA��9%����ҍ׾�H���z����F����/�`   `   hz̽L߽M�,I=�7�;w��4��2����7���W��tq��2��'���2���tq���W���7�2��4��;w��7�,I=�M�L߽`   `   43ٽZ��)��?�\����cؾ�?��;�ye��+���>���:���0���:���>���+��ye��;��?�cؾ���>�\�)��Z��`   `   ����D���9��%���&��z��2� �e��`��;N���r��)�Ϳ��Կ)�Ϳ�r��;N���`�� �e��2�z��&���%����9�D�`   `   �����&�X!]�K�����4��ZV�z���-����Ϳg#��£	�ɭ�£	�g#����Ϳ�-��z���ZV�4���K���X!]���&�`   `   ��0�<XE�e끾�_���w���9�x�x�֖��!:˿G���!�\;�\(E�\;���!�G�!:˿֖��w�x���9��w��_��e끾<XE�`   `   5O���e��~��@eҾ����R�^⋿tG��s��N#��Q���u��߁���u��Q�N#�s��tG��]⋿�R����@eҾ�~����e�`   `   �ln��#��������D�%�%�e�����09˿�
��DD����Ж��q���Ж����DD��
�09˿����%�e�D�%��������#��`   `   ����>���������1�us�䆡���ڿ��H�\�ԝ��g˪� ���g˪�ԝ��H�\�����ڿ䆡�us��1��������>��`   `   ����L��LȾv?���7��y��K��	῾�!�u�e�{Ж�,���@��,��{Ж�u�e���!�	��K���y���7�v?�LȾL��`   `   `,��J߳���վ�	�ԃ9�v�x�"q���3ܿ��?G]��ΐ�Vت����Vت��ΐ�?G]����3ܿ"q��v�x�ԃ9��	���վJ߳�`   `   ������ž���K\�r#7��oq��}����Ϳ��l'E����_Ж��R��_Ж����l'E�����Ϳ�}���oq�r#7�K\������ž`   `   d�Ѿ��ؾ���_�GF1��Ed�/��������)��D,$���Q��u�ו���u���Q�D,$��)������/����Ed�GF1��_��ﾠ�ؾ`   `   =��\1�f%��8C�?�(��R��%���-����Ϳ��[�!�q�:��DD�q�:�[�!�����Ϳ�-���%���R�?�(�8C�f%��\1�`   `   �Y��u�������'����K>�/�i��d�� ʫ��^ο,q�P�����P��,q��^ο ʫ��d��/�i�K>�����'����u���`   `   ^���)�u���	�D���(�I�<uq�U����O��غ��<˿B{ѿ�<˿غ��O��U���<uq�I���(�D��	�u���)�`   `   +��I��k������"�v2)���F�0�h�3ℿ6��w���w6��3ℿ0�h���F�v2)�"������k�I��`   `   ��$�)*�~� �F+��S� ��b������7�W}P�8�e���s���x���s�8�e�W}P���7�����b�S� �F+��~� �)*�$�`   `   d����
��{�������w�������-����p�,��:7��:��:7�p�,�����-�������w��徦���{���
�`   `   �E
�K*�^���=��hӾ��ž����L(Ⱦ��־;��N�����s����N���;�龲�־L(Ⱦ������žhӾ=��^���K*�`   `   ����|�ܢ��s�߾�nǾ1E��`���#-��7줾�0�����J^��2ڽ�J^������0��7줾#-��`���1E���nǾs�߾ܢ���|�`   `   �	�ƛ�s*������ž�ޫ������0��N5��{-��|��������4������|���{-��N5���0�������ޫ��ž���s*��ƛ�`   `   ��a�������Ҿl ��}�����KL`��L���@��6;�;�9��6;���@��L�KL`����}��l ���Ҿ�򾟨�a�`   `   x�,��(��g�a�����"ȾǢ��0��	�T�
1�h���W��#��W�h��
1�	�T��0��Ǣ��"Ⱦ���a��g��(�`   `   5�S�O�� A���+�b���@�8���������a�e-�\�	�g��J�۽g��\�	�e-���a�����8����@�b����+�� A�O�`   `   '���2���tq���W���7�2��4��;w��7�,I=�M�L߽hz̽L߽M�,I=�7�;w��4��2����7���W��tq��2��`   `   �0���:���>���+��ye��;��?�cؾ���?�\�)��Z��43ٽZ��)��?�\����cؾ�?��;�ye��+���>���:��`   `   ��Կ)�Ϳ�r��;N���`�� �e��2�z��&���%����9�D�����D���9��%���&��z��2� �e��`��;N���r��)�Ϳ`   `   ɭ�£	�g#����Ϳ�-��z���ZV�4���K���X!]���&������&�X!]�K�����4��ZV�z���-����Ϳg#��£	�`   `   \(E�\;���!�G�!:˿֖��w�x���9��w��_��e끾<XE���0�<XE�e끾�_���w���9�w�x�֖��!:˿G���!�\;�`   `   �߁���u��Q�N#�s��tG��]⋿�R����@eҾ�~����e�5O���e��~��@eҾ����R�]⋿tG��s��N#��Q���u�`   `   �q���Ж����DD��
�09˿����%�e�D�%��������#���ln��#��������D�%�%�e�����09˿�
��DD����Ж�`   `    ���g˪�ԝ��H�\�����ڿ䆡�us��1��������>������>���������1�us�䆡���ڿ��H�\�ԝ��g˪�`   `   �@��,��{Ж�u�e���!�	��K���y���7�v?�LȾL������L��LȾv?���7��y��K��	῾�!�u�e�{Ж�,��`   `   ���Vت��ΐ�?G]����3ܿ"q��v�x�ԃ9��	���վJ߳�`,��J߳���վ�	�ԃ9�v�x�"q���3ܿ��?G]��ΐ�Vت�`   `   �R��_Ж����l'E�����Ϳ�}���oq�r#7�K\������ž������ž���K\�r#7��oq��}����Ϳ��l'E����_Ж�`   `   ו���u���Q�D,$��)������/����Ed�GF1��_��ﾠ�ؾd�Ѿ��ؾ���_�GF1��Ed�/��������)��D,$���Q��u�`   `   �DD�q�:�[�!�����Ϳ�-���%���R�?�(�8C�f%��\1�=��\1�f%��8C�?�(��R��%���-����Ϳ��[�!�q�:�`   `   ���P��,q��^ο ʫ��d��/�i�K>�����'����u����Y��u�������'����K>�/�i��d�� ʫ��^ο,q�P��`   `   C{ѿ�<˿غ��O��U���<uq�I���(�D��	�u���)�^���)�u���	�D���(�I�<uq�U����O��غ��<˿`   `   ���w6��3ℿ0�h���F�v2)�"������k�I��+��I��k������"�v2)���F�0�h�3ℿ6��w`   `   ��x���s�8�e�W}P���7�����b�S� �F+��~� �)*�$���$�)*�~� �F+��S� ��b������7�W}P�8�e���s�`   `   �:��:7�p�,�����-�������w��徦���{���
�d����
��{�������w�������-����p�,��:7�`   `   s����N���;�龲�־L(Ⱦ������žhӾ=��^���K*��E
�K*�^���=��hӾ��ž����L(Ⱦ��־;��N�����`   `   2ڽ�J^������0��7줾#-��`���1E���nǾs�߾ܢ���|�����|�ܢ��s�߾�nǾ1E��`���#-��7줾�0�����J^��`   `   �4������|���{-��O5���0�������ޫ��ž���s*��Ǜ��	�Ǜ�s*������ž�ޫ������0��N5��{-��|�������`   `   ;�9��6;���@��L�KL`����}��l ���Ҿ�򾟨�a���a�������Ҿl ��}�����KL`��L���@��6;�`   `   �#��W�h��
1�	�T��0��Ǣ��"Ⱦ���a��g��(�x�,��(��g�a�����"ȾǢ��0��	�T�
1�h���W�`   `   J�۽g��\�	�e-���a�����8����@�b����+�� A�O�5�S�O�� A���+�b���@�8���������a�e-�\�	�g��`   `   =������&�M���[����8ƾ4���W��Q�7��N���]�c���]��N�Q�7�W��4���8ƾ����[�M���&����`   `   �f����ƽ3����7�T���Q��z��oW���=��_��y�Z�������Z����y��_���=�nW�z��Q��T�����7�3����ƽ`   `   "Gнl�MA�L�Z�����ؾ��t�;��f��c���d���R��UD���R���d���c���f�t�;����ؾ���L�Z�MA�l�`   `   I��i���8�D��3]���G�%.�uB_�<��pȟ�?.���ſ�
˿�ſ?.��pȟ�<��uB_�%.��G�3]��D���8�i��`   `   �;�ߑ)�ߏ[������ؾu��;J�������������0�ۿ����Ud������0�ۿ������������;J�u����ؾ���ߏ[�ߑ)�`   `   ��8��vJ��s��������=�*���c���������6ݿ�,��������,�6ݿ����������c�=�*��������s���vJ�`   `   ��\�!$o�	퓾=ƾ���0�;��x�!���_nǿ���"~���4�0�=���4�"~����_nǿ!����x�0�;����=ƾ	퓾!$o�`   `   o_���S��AQ����ھ����G�]��V���ֿ�
���-��J��T��J���-��
��ֿV��]����G�����ھAQ���S��`   `   Ep��+���UX�����y��O�\b���媿K�ۿ�^�s�4�JR�VJ]�JR�s�4��^�K�ۿ�媿\b��O�y�����UX��+���`   `   �������,׾q" ��!��%Q�l酿�Ȩ��:׿��{4.��#J���T��#J�{4.����:׿�Ȩ�l酿�%Q��!�q" ��,׾���`   `   f�ྵ����ՠ	�� %�ĞN�䁿�Q���ɿ:c�����f�4�Y�=�f�4����:c���ɿ�Q��䁿ĞN�� %�ՠ	�����`   `   Ao����e
�]���J'��UH���u��蕿Xc����޿:e��W��E��W�:e���޿Xc���蕿��u��UH��J'�]���e
���`   `   g�L �mV��$��u(��K?�<c��⇿�R��l����ۿ����������ۿl���R���⇿<c��K?��u(��$�mV�L �`   `   m 8�=5�(.��(�Ϛ(��s4�?M�/p�$���à�j��Aÿi�ȿAÿj���à�$��/p�?M��s4�Ϛ(��(�(.�=5�`   `   #�M��*I�0V=�i�/�b,'��w(��6��N��dm��e��#.���㝿(o���㝿#.���e���dm��N��6��w(�b,'�i�/�0V=��*I�`   `   1�\���V��G�ɕ3�dN#�����0�.~-�� C�z�Z�>�o��6~�����6~�>�o�z�Z�� C�.~-��0����dN#�ɕ3��G���V�`   `   $b�(J[�d+I���1�Y�y� �	�U����.B,�G�;�8jF�eDJ�8jF�G�;�.B,����U� �	�y�Y���1�d+I�(J[�`   `   L]��V�6LC��*��d�@ ��B����������9��f~�9����������龁B�@ ��d��*�6LC��V�`   `   ��O�+I��=7���y�����YeʾLi���y���(ƾ7hо�ؾ��۾�ؾ7hо�(ƾ�y��Li��Yeʾ���y�����=7�+I�`   `   W�>���8�Ͳ(��n����@S;�2��~z��^Y��Q������A ������Q��^Y��z��~�2��@S;����n�Ͳ(���8�`   `   _�/���*�\X��C�2��gż�~������Fo��a���[�+�Z�!�Z�+�Z���[��a�Fo�����~��gż�2�侢C�\X���*�`   `   �Y(�0�#�)���H���޾Bɶ�r-�� -r��jK�,2��c#�����������c#�,2��jK� -r�r-��Bɶ���޾�H�)��0�#�`   `   �,�.w(�����	����9d���՗�>o�D=��Q���^8齻��^8����Q�D=�>o��՗�9d������	����.w(�`   `   �}@���;��n.�C����D�վ1o���G��VWC�T���|��������������|�T��VWC��G��1o��D�վ��C���n.���;�`   `   c���]��N�Q�7�W��4���8ƾ����[�M���&����=������&�M���[����8ƾ4���W��Q�7��N���]�`   `   ����Z����y��_���=�nW�z��Q��T�����7�3����ƽ�f����ƽ3����7�T���Q��z��nW���=��_��y�Z���`   `   UD���R���d���c���f�t�;����ؾ���L�Z�MA�l�#Gнl�MA�L�Z�����ؾ��t�;��f��c���d���R��`   `   �
˿�ſ?.��pȟ�<��uB_�%.��G�3]��D���8�j��J��j���8�D��3]���G�%.�uB_�<��pȟ�?.���ſ`   `   Ud������0�ۿ������������;J�u����ؾ���ߏ[�ߑ)��;�ߑ)�ߏ[������ؾu��;J�������������0�ۿ����`   `   �����,�6ݿ����������c�=�*��������s���vJ���8��vJ��s��������=�*���c���������6ݿ�,���`   `   0�=���4�"~����_nǿ!����x�0�;����=ƾ	퓾!$o���\�!$o�	퓾=ƾ���0�;��x�!���_nǿ���"~���4�`   `   �T��J���-��
��ֿV��]����G�����ھAQ���S��o_���S��AQ����ھ����G�]��V���ֿ�
���-��J�`   `   VJ]�JR�s�4��^�K�ۿ�媿\b��O�y�����UX��+���Ep��+���UX�����y��O�\b���媿K�ۿ�^�s�4�JR�`   `   ��T��#J�{4.����:׿�Ȩ�l酿�%Q��!�q" ��,׾����������,׾q" ��!��%Q�l酿�Ȩ��:׿��{4.��#J�`   `   Y�=�f�4����:c���ɿ�Q��䁿ĞN�� %�ՠ	�����f�ྵ����ՠ	�� %�ĞN�䁿�Q���ɿ:c�����f�4�`   `   �E��W�:e���޿Xc���蕿��u��UH��J'�]���e
���Ao����e
�]���J'��UH���u��蕿Xc����޿:e��W�`   `   �������ۿl���R���⇿<c��K?��u(��$�mV�L �g�L �mV��$��u(��K?�<c��⇿�R��l����ۿ���`   `   i�ȿAÿj���à�$��/p�?M��s4�Ϛ(��(�(.�=5�m 8�=5�(.��(�Ϛ(��s4�?M�/p�$���à�j��Aÿ`   `   (o���㝿#.���e���dm��N��6��w(�c,'�i�/�0V=��*I�#�M��*I�0V=�i�/�b,'��w(��6��N��dm��e��#.���㝿`   `   ����6~�>�o�z�Z�� C�.~-��0����dN#�ɕ3��G���V�1�\���V��G�ɕ3�dN#�����0�.~-�� C�z�Z�>�o��6~�`   `   eDJ�8jF�G�;�.B,����U� �	�y�Y���1�d+I�(J[�$b�(J[�d+I���1�Y�y� �	�U����.B,�G�;�8jF�`   `   f~�9����������龁B�@ ��d��*�6LC��V�L]��V�6LC��*��d�@ ��B����������9��`   `   ��۾�ؾ7hо�(ƾ�y��Li��Yeʾ���y�����=7�+I���O�+I��=7���y�����YeʾLi���y���(ƾ7hо�ؾ`   `   A ������Q��^Y��z��~�2��@S;����n�Ͳ(���8�W�>���8�Ͳ(��n����@S;�2��}z��^Y��Q������`   `   !�Z�+�Z���[��a�Fo�����~��gż�2�侢C�\X���*�_�/���*�\X��C�2��gż�~������Fo��a���[�+�Z�`   `   �������c#�,2��jK�!-r�r-��Bɶ���޾�H�)��0�#��Y(�0�#�)���H���޾Bɶ�r-�� -r��jK�,2��c#����`   `   ���^8����Q�D=�>o��՗�9d������	����.w(��,�.w(�����	����9d���՗�>o�D=��Q���^8�`   `   ���������|�T��VWC��G��1o��D�վ��C���n.���;��}@���;��n.�C����D�վ1o���G��VWC�T���|�����`   `   &���cȑ�&���,���7��n|��G��@Xؾ��w3���2�ڬ@�g�E�ڬ@���2�w3���@Xؾ�G���n|��7�,��&���cȑ�`   `   憍��z��J�ѽm����R�<đ���¾%,�����5�oBL�)[�\[`�)[�oBL��5���%,����¾<đ���R�m��I�ѽ�z��`   `   R������������/��x�����澂����5��GU�Ʊn�_8��{��_8�Ʊn��GU���5����������x���/��������`   `   w�ҽ.L齈���Q�	7����ʾ���b	.��1U� �x��׊��n��K՗��n���׊� �x��1U�b	.������ʾ	7����Q���.L�`   `   �.�6��~7���x����l�뾙��C�H���t��o��~���u�����u���~����o����t�C�H����l�뾄����x�~7�6��`   `   ��(�r�5�Gu]�6����Už����0��`����������Ǵ�q�ĿZyʿq�Ŀ�Ǵ����������`���0����Už6���Gu]�r�5�`   `   �U�Mb���?����ݾ�����A�C�t��<��B����zȿQ}ܿ�/�Q}ܿ�zȿB����<��C�t���A������ݾ?����Mb�`   `   ��	���f���@���k����n�<N�x����B���w����ֿ�n�$����n�ֿ�w���B��x���<N��n�k���@���f���	���`   `   �Ԯ����\���ܾA���@(��EU��$�� ���횽�	}ܿk,������k,��	}ܿ횽� ����$���EU��@(�A���ܾ\�����`   `   ?��Fk�>������l�.�@XW�֘�� ���;'��J׿3�Y|��3�J׿;'�� ���֘��@XW�l�.����>���Fk��`   `   �����������@�2���T��7����������ȿO}ܿ`�O}ܿ��ȿ��������7���T�@�2���������`   `   @<���8��V1��*��m*�@�5�]�N��gq�����ra��A2��+;Ŀ��ɿ+;ĿA2��ra�������gq�]�N�@�5��m*��*��V1���8�`   `   �2l��0f��V��0E���8�*,8��E�
_��9��U������K���о��K��������U���9�
_��E�*,8���8��0E��V��0f�`   `   �j���؊�o�}��g`��G��s9���:��I�mua�^�{�N���B�����B��N���^�{�mua��I���:��s9��G��g`�o�}��؊�`   `   �h��SV���d���'x�ЯR���8��.���2�i�A�LU�5�g�ʚt�:y�ʚt�5�g�LU�i�A���2��.���8�ЯR��'x��d��SV��`   `   ���|��Fq���؃���X�TG5�rF!�R1�y"��.�JE<�pF��I�pF�JE<��.�y"�R1�rF!�TG5���X��؃�Fq��|��`   `   �����ڴ�uV��ϓ��y�V��y-�������F��%������z�����z����%��F���������y-�y�V�ϓ��uV���ڴ�`   `   �ɶ��:��� ��'����L�#F!�bR�!)���ؾ�\ھ�
⾉y��p쾉y龖
��\ھ��ؾ!)�bR�#F!��L�'���� ���:��`   `   ���1V���>���4l� 7;���������s8��oP���N���!���u���!���N��oP��s8���������� 7;��4l��>��1V��`   `   Kԑ��2���z���P��-&�f� ���Ⱦ1��𙋾U�.�y�Z�x���x�Z�x�.�y�U�𙋾1����Ⱦf� ��-&���P��z��2��`   `   %'x�:9o�B�V��b5�	�����ᮾ�����jb�5F���7��`1��/��`1���7�5F��jb������ᮾ��	���b5�B�V�:9o�`   `   tT�|M�?P:��S�N����˾�Ꜿ�q���>����	�����x��������	�����>��q��Ꜿ��˾N���S�?P:�|M�`   `   p�>�K�8�VH)�2��.��I�� ��Ddb�{�+�&B�!rؽ�����᳽����!rؽ&B�{�+�Ddb� ��I��.��2��VH)�K�8�`   `   �k9�c{4�V�&�p8����x�ľ_Ř��f�^�)��C��c���]�������]��c���C��^�)��f�_Ř�x�ľ���p8�V�&�c{4�`   `   g�E�ڬ@���2�w3���@Xؾ�G���n|��7�,��&���dȑ�&���dȑ�&���,���7��n|��G��@Xؾ��w3���2�ڬ@�`   `   \[`�)[�oBL��5���%,����¾<đ���R�m��J�ѽ�z��憍��z��J�ѽm����R�<đ���¾%,�����5�oBL�)[�`   `   �{��_8�Ʊn��GU���5����������x���/��������R������������/��x�����澁����5��GU�Ʊn�_8�`   `   K՗��n���׊� �x��1U�b	.������ʾ	7����Q���.L�w�ҽ.L齈���Q�	7����ʾ���b	.��1U� �x��׊��n��`   `   ��u���~����o����t�C�H����l�뾄����x�~7�6���.�6��~7���x����l�뾙��C�H���t��o��~���u���`   `   Zyʿq�Ŀ�Ǵ����������`���0����Už6���Gu]�r�5���(�r�5�Gu]�6����Už����0��`����������Ǵ�q�Ŀ`   `   �/�Q}ܿ�zȿB����<��C�t���A������ݾ?����Mb��U�Mb���?����ݾ�����A�C�t��<��B����zȿQ}ܿ`   `   $����n�ֿ�w���B��x���<N��n�k���@���f���	�����	���f���@���k����n�<N�x����B���w����ֿ�n�`   `   ����k,��	}ܿ횽� ����$���EU��@(�A���ܾ\������Ԯ����\���ܾA���@(��EU��$�� ���횽�	}ܿk,��`   `   Y|��3�J׿;'�� ���֘��@XW�l�.����>���Fk��?��Fk�>������l�.�@XW�֘�� ���;'��J׿3�`   `   `�O}ܿ��ȿ��������7���T�@�2��������������������@�2���T��7����������ȿO}ܿ`   `   ��ɿ+;ĿA2��ra�������gq�]�N�@�5��m*��*��V1���8�@<���8��V1��*��m*�@�5�]�N��gq�����ra��A2��+;Ŀ`   `   о��K��������U���9�
_��E�*,8���8��0E��V��0f��2l��0f��V��0E���8�*,8��E�
_��9��U������K���`   `   ���B��N���^�{�mua��I���:��s9��G��g`�o�}��؊��j���؊�o�}��g`��G��s9���:��I�mua�^�{�N���B��`   `   :y�ʚt�5�g�LU�i�A���2��.���8�ЯR��'x��d��SV���h��SV���d���'x�ЯR���8��.���2�i�A�LU�5�g�ʚt�`   `   �I�pF�JE<��.�y"�R1�rF!�TG5���X��؃�Fq��|�����|��Fq���؃���X�TG5�rF!�R1�y"��.�JE<�pF�`   `   ����z����%��F���������y-�y�V�ϓ��uV���ڴ������ڴ�uV��ϓ��y�V��y-�������F��%������z�`   `   �p쾉y龖
��\ھ��ؾ!)�bR�$F!��L�'���� ���:���ɶ��:��� ��'����L�#F!�bR�!)���ؾ�\ھ�
⾉y�`   `   �u���!���N��oP��s8���������� 7;��4l��>��1V�����1V���>���4l� 7;���������s8��oP���N���!��`   `   ��x�Z�x�.�y�U�𙋾1����Ⱦf� ��-&���P��z��2��Kԑ��2���z���P��-&�f� ���Ⱦ1��𙋾U�.�y�Z�x�`   `   �/��`1���7�5F��jb������ᮾ��	���b5�B�V�:9o�%'x�:9o�B�V��b5�	�����ᮾ�����jb�4F���7��`1�`   `   x��������	�����>��q��Ꜿ��˾N���S�?P:�|M�tT�|M�?P:��S�N����˾�Ꜿ�q���>����	�����`   `   �᳽����!rؽ&B�{�+�Ddb� ��I��.��2��VH)�K�8�p�>�K�8�UH)�1��.��I�� ��Ddb�{�+�&B�!rؽ����`   `   �����]��c���C��_�)��f�_Ř�x�ľ���p8�V�&�c{4��k9�c{4�V�&�p8����x�ľ_Ř��f�^�)��C��c���]��`   `   ,�I�׀b�8���K�׽s��Y������r��/U�;� %#���0�f�5���0� %#�;�/Uﾨr������Y�s��K�׽7���׀b�`   `   [��Rw��֥�J���)�
ul������0̾fG���*��s(��T5���9��T5��s(��*�fG���0̾����
ul���)�I���֥��Rw�`   `   Az��>�i�Ž��
���C�ͅ���겾��6���]%�r�9��)G�	�K��)G�r�9��]%�6�����겾ͅ����C���
�i�Ž>�`   `   ������½ ���!�&�)De�3����|;3��ph �v�;��5R�O�`�,�e�O�`��5R�v�;�ph �3���|;3���(De�!�&� �����½`   `   �f�����G��FII�˂��ׇ��
 뾓K�o46�8�T��l���|������|��l�8�T�o46��K�
 �ׇ��˂��FII�G������`   `   /]!���)��WD��"s�����Yo̾�V��	'���J���k�|��ֶ���Ŏ�ֶ��|����k���J��	'��V�Yo̾�����"s��WD���)�`   `   �"\��kc�.�z��쒾ϴ���侚���36���[��x~��f�������f�������f���x~���[��36�������ϴ��쒾.�z��kc�`   `   X���-љ�ۡ�Й����Ͼ������DbA���g�A���5b�� ���
f�� ���5b��A�����g�DbA���������ϾЙ��ۡ�-љ�`   `   2<Ҿ�(Ҿ7�Ӿ��۾�Nﾪ�	�r\%���G��l�#�������r���F���r������#���l���G�r\%���	��Nﾯ�۾7�Ӿ�(Ҿ`   `   �?��O��������
�	��s~+��I���k��w��6��������`������6����w����k��I�s~+�	����
�������O�`   `   gFJ��E��m9���+�Uy"��$#���/�,*G�wd� ��$ ��X���e:��X���$ �� ��wd�,*G���/��$#�Uy"���+��m9��E�`   `   픉��6��l�s�SrW��6?�i2�13��4A�I�W���p�힃��U��D���U��힃���p�I�W��4A�13�i2��6?�SrW�l�s��6��`   `   �赿b﮿J����t���!`�wfB�?�5���8�",G�B�Z���l� �y��{~� �y���l�A�Z�",G���8�?�5�wfB��!`��t��J���b﮿`   `   W��ϼܿ�a¿ˠ�b"��7�R�c57��.�P�3��@�v�N��Y���\��Y�v�N��@�P�3��.�c57�7�R�b"��ˠ��a¿ϼܿ`   `   g�
�������Ź��B��a#`�:�6�N(#�^w��a%���.�t96�9�t96���.��a%�^w�N(#�:�6�a#`��B���Ź���忍�`   `   @��?�����eX˿�Q���eg��3�C���+��
��1�����������1��
��+�C���3��eg��Q��eX˿���?��`   `   �3"�M�����ѿH���äe���+�t��R\��5�(	�-��,�-�(	��5�R\�t����+�äe�H����ѿ��M��`   `   ���\���2��4Kɿ�P����Y�W��u�ʹʾ�����F���8�������8���F������ʹʾu�W����Y��P��4Kɿ�2��\��`   `   #�
�Y�Q:�'鵿Kw����E�A�\�Ӿ�������ę��������ę���������\�ӾA���E�Kw��'鵿Q:�Y�`   `   �S�C�ݿJ"��챛�|*l��	,�
��Qz�������g���O�ƕE���B�ƕE���O��g�����Qz��
���	,�|*l�챛�J"��C�ݿ`   `   gŹ��ݱ�v���&-����E����
HҾI��i�c���4�����t�+�
��t������4�i�c�I��
HҾ�����E�&-��v����ݱ�`   `   ����!����y�U�O��S#�qu��(���8����<�A������̽o�ý��̽��A����<��8��(��qu���S#�U�O���y�!��`   `   zh�#!`��NJ��+���	���Ӿ��#�c�ʌ#����s������3�����s�����ʌ#�#�c�����Ӿ��	��+��NJ�#!`�`   `   
�C�� >��-���6v������P'��W�U�DU��Q׽����Zs�]�Zs������Q׽DU�W�U�P'������6v�����-�� >�`   `   f�5���0� %#�;�/Uﾨr������Y�s��K�׽8���׀b�,�I�׀b�8���K�׽s��Y������r��/U�;� %#���0�`   `   ��9��T5��s(��*�fG���0̾����
ul���)�J���֥��Rw�[��Rw��֥�J���)�
ul������0̾fG���*��s(��T5�`   `   �K��)G�r�9��]%�6�����겾ͅ����C���
�i�Ž>�Az��>�i�Ž��
���C�ͅ���겾��6���]%�r�9��)G�`   `   ,�e�O�`��5R�v�;�ph �3���|;3���)De�!�&� �����½������½ ���!�&�)De�3����|;3��ph �v�;��5R�O�`�`   `   �����|��l�8�T�o46��K�
 �ׇ��˂��FII�G�������f�����G��FII�˂��ׇ��
 뾓K�o46�8�T��l���|�`   `   �Ŏ�ֶ��|����k���J��	'��V�Yo̾�����"s��WD���)�/]!���)��WD��"s�����Yo̾�V��	'���J���k�|��ֶ��`   `   �f�������f���x~���[��36�������ϴ��쒾.�z��kc��"\��kc�.�z��쒾ϴ���侚���36���[��x~��f������`   `   
f�� ���5b��A�����g�DbA���������ϾЙ��ۡ�-љ�X���-љ�ۡ�Й����Ͼ������DbA���g�A���5b�� ���`   `   �F���r������#���l���G�r\%���	��Nﾯ�۾7�Ӿ�(Ҿ2<Ҿ�(Ҿ7�Ӿ��۾�Nﾪ�	�r\%���G��l�#�������r��`   `   �`������6����w����k��I�s~+�	����
�������O��?��O��������
�	��s~+��I���k��w��6�������`   `   e:��X���$ �� ��wd�,*G���/��$#�Uy"���+��m9��E�gFJ��E��m9���+�Uy"��$#���/�,*G�wd� ��$ ��X���`   `   D���U��힃���p�I�W��4A�13�i2��6?�SrW�l�s��6��픉��6��l�s�SrW��6?�i2�13��4A�I�W���p�힃��U��`   `   �{~� �y���l�B�Z�",G���8�?�5�wfB��!`��t��J���b﮿�赿b﮿J����t���!`�wfB�?�5���8�",G�B�Z���l� �y�`   `   ��\��Y�v�N��@�P�3��.�c57�7�R�b"��ˠ��a¿ϼܿW��ϼܿ�a¿ˠ�b"��7�R�c57��.�P�3��@�v�N��Y�`   `   9�t96���.��a%�^w�N(#�:�6�a#`��B���Ź���忍�g�
�������Ź��B��a#`�:�6�N(#�^w��a%���.�t96�`   `   �������1��
��+�C���3��eg��Q��eX˿���?��@��?�����eX˿�Q���eg��3�C���+��
��1����`   `   �,�-�(	��5�R\�t����+�äe�H����ѿ��M���3"�M�����ѿG���äe���+�t��R\��5�(	�-�`   `   �����8���F������ʹʾu�W����Y��P��4Kɿ�2��\�����\���2��4Kɿ�P����Y�W��u�ʹʾ�����F���8��`   `   �����ę���������\�ӾA���E�Kw��'鵿Q:�Y�#�
�Y�Q:�'鵿Kw����E�A�\�Ӿ�������ę���`   `   ��B�ƕE���O��g�����Qz��
���	,�|*l�챛�J"��C�ݿ�S�C�ݿJ"��챛�{*l��	,�
��Qz�������g���O�ƕE�`   `   +�
��t������4�i�c�I��
HҾ�����E�&-��v����ݱ�gŹ��ݱ�v���&-����E����
HҾI��i�c���4�����t�`   `   o�ý��̽��A����<��8��(��qu���S#�V�O���y�!������!����y�U�O��S#�qu��(���8����<�A������̽`   `   �3�����s�����ʌ#�#�c�����Ӿ��	��+��NJ�#!`�zh�#!`��NJ��+���	���Ӿ��#�c�ʌ#����s�����`   `   ]�Zs������Q׽DU�W�U�P'������7v�����-�� >�
�C�� >��-���6v������P'��W�U�DU��Q׽����Zs�`   `   ,��
0��t�&�����B�����e���[%従^��
!�� 0�B]5�� 0��
!��^�[%�e��������B���&���t�
0�`   `   OM*��:A�����ZT��<�
��vC��|��c����־l& �[����h�!���[��l& ���־c���|���vC�<�
�ZT�������:A�`   `   �1]�C�t�B4���O۽l��dR�����ݛ��@n۾�+�h��9�� ��9�h��+�@n۾ݛ�������dR�l��O۽B4��C�t�`   `   
S���&���O˽����1��ql�����by¾���|
����&���)��&���|
����by¾�����ql���1����O˽�&��`   `   �����&��h%��_R��a��Yݬ�P�׾����B��*���5���9���5��*��B����P�׾Yݬ��a���_R��h%�&���`   `   ��#��t(�U�6���Q�~�{��������QHﾐ���'�:��rF���J��rF�:��'����QHﾛ������~�{���Q�U�6��t(�`   `   Q�p�F#s�$`{�s���嗾�����׾*�����O�3�X�G���T��IY���T�X�G�O�3����*���׾����嗾s���$`{�F#s�`   `   ޱ��ٰ�c2������9����̾�	����$�m	=��&Q�F[^���b�F[^��&Q�m	=���$���	��̾�9�����c2���ٰ�`   `   h���;������꾾徚�+�P^�B*�\.A��T�u�a�LXf�u�a��T�\.A�B*�P^�+��쾾��꾗����;�`   `   +�A��<�_�.�x�����/0	�9E���O+��@�;R�	�^�{�b�	�^�;R��@�O+���9E�/0	����x��_�.��<�`   `   (W��{b��@�v�?GU�N\6��
!���:�V�(�\�9�v�I���T���X���T�u�I�\�9�V�(��:���
!�N\6�?GU�@�v�{b��`   `   eʿ�����]���Ǝ��9g�'>��J&���$�#�*4/�P�;��BE���H��BE�P�;�*4/�$�#����J&�'>��9g��Ǝ��]������`   `   
M�ނ�1��(���Ǜ����_��_5�:� �x<��j!�{
*��91���3��91�{
*��j!�x<�:� ��_5���_�Ǜ��(���1��ނ�`   `   �:��{0��X��������z(���VD���!��c��������e�GM��e��������c���!��VD�z(����������X��{0�`   `   �>j��\��e8��Z��̿U���|�P��!�	�/��� ���r������ �/�	��!�|�P�U����̿�Z��e8��\�`   `   ���2~�[NR����s�࿋뚿�(W�����0���s�/�ؾ�׾ؾ�׾/�ؾ�s��0������(W��뚿s�࿾��[NR�2~�`   `   B2��蛅��\��$�۴翮W��KU�?5��*�ߒ������Э�>嬾�Э����ߒ���*�?5�KU��W��۴��$��\�蛅�`   `   ���R~�<R�����޿ʖ�g
J�>�
�W�ʾ'C���n��߈�����߈��n��'C��W�ʾ>�
�g
J�ʖ���޿��<R�R~�`   `   �Vj�I\�-8�M���ǿ<d����6������A��"����d��nR�C_M��nR��d�"����A��������6�<d����ǿM�-8�I\�`   `   �;�
�0��D�����j����*wԾ����"�Z��`1��������`1�"�Z�����*wԾ����j����D��
�0�`   `   VZ��Q���1ѷ��c��&�@�v��ȡ��P7s�|_.�� �r�D_۽r罴 �|_.�P7s�ȡ��v��&�@��c��1ѷ����Q�`   `   �ο:�ſ�,���n��{�U�[S�]�־�Z��l�F�T|
��̽�����f�������̽T|
�l�F��Z��]�־[S�{�U��n���,��:�ſ`   `   ��� ���~���	IU�}r&�x�����65s� %����[V����t��2^���t�[V����� %�65s���x���}r&�	IU�~��� ���`   `   �~a�-�Y���D�h�&�S��s�˾.��y0R����x���2��V�@��*�V�@�2��x������y0R�.��s�˾S��h�&���D�-�Y�`   `   B]5�� 0��
!��^�[%�e��������B���&���t�
0�,��
0��t�&�����B�����e���[%従^��
!�� 0�`   `   h�!���[��l& ���־c���|���vC�<�
�ZT�������:A�PM*��:A�����ZT��<�
��vC��|��c����־l& �[����`   `   � ��9�h��+�@n۾ݛ�������dR�l��O۽B4��C�t��1]�C�t�B4���O۽l��dR�����ݛ��@n۾�+�h��9�`   `   ��)��&���|
����by¾�����ql���1����O˽�&��S���&���O˽����1��ql�����by¾���|
����&�`   `   ��9���5��*��B����P�׾Yݬ��a���_R��h%�&��������&��h%��_R��a��Yݬ�P�׾����B��*���5�`   `   ��J��rF�:��'����QHﾛ������~�{���Q�U�6��t(���#��t(�U�6���Q�~�{��������QHﾐ���'�:��rF�`   `   �IY���T�X�G�O�3����*���׾����嗾s���$`{�F#s�Q�p�F#s�$`{�s���嗾�����׾*�����O�3�X�G���T�`   `   ��b�F[^��&Q�m	=���$���	��̾�9�����c2���ٰ�ޱ��ٰ�c2������9����̾�	����$�m	=��&Q�F[^�`   `   LXf�u�a��T�\.A�B*�P^�+��쾾��꾗����;�h���;������꾾徚�+�P^�B*�\.A��T�u�a�`   `   {�b�	�^�;R��@�O+���9E�/0	����x��_�.��<�+�A��<�_�.�x�����/0	�9E���O+��@�;R�	�^�`   `   ��X���T�v�I�\�9�V�(��:���
!�N\6�?GU�@�v�{b��(W��{b��@�v�?GU�N\6��
!���:�V�(�\�9�v�I���T�`   `   ��H��BE�P�;�*4/�$�#����J&�'>��9g��Ǝ��]������eʿ�����]���Ǝ��9g�'>��J&���$�#�*4/�P�;��BE�`   `   ��3��91�{
*��j!�x<�:� ��_5���_�Ǜ��(���1��ނ�
M�ނ�1��(���Ǜ����_��_5�:� �x<��j!�{
*��91�`   `   GM��e��������c���!��VD�z(����������X��{0��:��{0��X��������z(���VD���!��c��������e�`   `   r������ �/�	��!�|�P�U����̿�Z��e8��\��>j��\��e8��Z��̿U���|�P��!�	�/��� ���`   `   ؾ�׾/�ؾ�s��0������(W��뚿s�࿾��[NR�2~����2~�[NR����s�࿋뚿�(W�����0���s�/�ؾ�׾`   `   >嬾�Э����ߒ���*�?5�KU��W��۴��$��\�蛅�B2��蛅��\��$�۴翮W��KU�?5��*�ߒ������Э�`   `   ����߈��n��'C��W�ʾ>�
�g
J�ʖ���޿��<R�R~����R~�<R�����޿ʖ�g
J�>�
�W�ʾ'C���n��߈�`   `   C_M��nR��d�"����A��������6�<d����ǿM�-8�I\��Vj�I\�-8�M���ǿ<d����6������A��"����d��nR�`   `   �����`1�"�Z�����*wԾ����j����D��
�0��;�
�0��D�����j����*wԾ����"�Z��`1���`   `   D_۽r罴 �|_.�P7s�ȡ��v��&�@��c��1ѷ����Q�VZ��Q���0ѷ��c��&�@�v��ȡ��P7s�|_.�� �r�`   `   �f�������̽T|
�m�F��Z��]�־[S�{�U��n���,��:�ſ�ο:�ſ�,���n��{�U�[S�]�־�Z��l�F�T|
��̽����`   `   �2^���t�[V����� %�65s���x���}r&�	IU�~��� ������ ���~���	IU�}r&�x�����65s� %����[V����t�`   `   �*�V�@�2��x������y0R�.��s�˾S��h�&���D�-�Y��~a�-�Y���D�h�&�S��s�˾.��y0R����x���2��V�@�`   `   �o��K���N��Ѡ������7���{��
���$:*��;�3SB��;�$:*��
��{������7�����Ѡ���N��K�`   `   �{�>���W�l䞽�`꽽�'���g��<��$¾���U��C��Z9�C��U�����$¾�<����g���'��`�l䞽�W�>��`   `   �<�+~N��R�����?@���'��;_��r���A����ѾQd�F����7�F���Qd��Ѿ�A���r���;_��'�?@������R��+~N�`   `   
<���󖽏ܮ���ؽ8m�z�4�� h��Z��{9����;H�[���)m��[���H澉�;{9���Z��� h�z�4�8m���ؽ�ܮ���`   `   ]?߽n��Cp������'��gM�y�}��������־�.�/G�����/G���.�־�������y�}��gM��'����Cp��n��`   `   ��.��/�_�3�)�=��,Q��bp�v���9����ƾt0侼���b��ߦ	�b������t0���ƾ9��v����bp��,Q�)�=�_�3��/�`   `   �N�����h������eㅾ�o������v��[�վ�"�o+�o��*��o��o+��"�[�վv�������o��eㅾ���h������`   `    7Ծо�8ž�s���;��&�����T�ɾ�h�T@�������������T@���h�T�ɾ���&���;���s���8žо`   `   Tz$�����d��t�:��E�־q�Ѿ}�ھx0�8������d�������8�x0�}�ھq�ѾE�־:���t��d����`   `   9}�Tt���[��_<����������R��B������g�����k����g�����B���R�쾏���������_<���[�Tt�`   `   K����c�������m��q�U��:*�������������9��X�����X��9���������������:*�q�U��m�������c��`   `   j;�!
	���쿉��֩��&AW��^&���
��,���x���#�|����|���#��x���,����
��^&�&AW�֩��������!
	�`   `   �S���F�R�'��|�찼��3���UB�/&�����D�ﾻ2�Md�8%�Md�2�D�ﾴ���/&��UB��3��찼��|�R�'���F�`   `   ㄕ��?��LYd�nG*�������!_��O!�[���!���a׾��վe�վ��վ�a׾!��[����O!��!_��������nG*�LYd��?��`   `   �?����������vS��f�����yx��<*��T����Ѿ�[�� ���ʷ� ���[����Ѿ�T���<*��yx�����f��vS��������`   `   N����������|s�J)!��)Ͽ;�����.�i]������k,������^������k,������i]����.�;����)ϿJ)!��|s��������`   `   *��A�����̾�f�'�uFտo����,�ӷ��v��Yt��p]���}�p]��Yt���v��ӷ龻�,�o��uFտf�'�̾����A��`   `   �������	��>Us��� �1ͿJ߀�2#�2�־DӘ��@q���S�CgK���S��@q�DӘ�2�־2#�J߀�1Ϳ�� �>Us��	������`   `   �?������ג��S��b�e���yi��h��þ�A��4*F���'�o����'�4*F�A���þ��h��yi�e���b��S��ג����`   `   ����E��l>d�Ǳ)��뿴 ��نH�F����C��a�Z�=��&;����&;�=��a�Z��C��F���نH�� ����Ǳ)�l>d��E��`   `   ?vS�4G��'�=� �e����z�h~$��*Ӿ�#��R.1�k}��Cz�����Cz��k}��R.1��#���*Ӿh~$���z�e��=� ��'�4G�`   `   G�v�	�"��ݻ�����(B��`�i�� AZ�9��w���z��b}��z��w��9�� AZ�i���`�(B�����ݻ�"��v�	�`   `   nWſ񯼿����Yn��]�L��h��;˾$����.�lO߽�/��ƅN��;4�ƅN��/��lO߽��.�$���;˾�h�^�L�Yn������񯼿`   `   L���wX����h�:�A�)���?��ҟ���Y�������">h�6�����6��">h���������Y��ҟ��?�)��:�A���h�wX��`   `   3SB��;�$:*��
��{������7�����Ѡ���N��K��o��K���N��Ѡ������7���{��
���$:*��;�`   `   Z9�C��U�����$¾�<����g���'��`�l䞽�W�>���{�>���W�l䞽�`꽽�'���g��<��$¾���U��C��`   `   �7�F���Qd��Ѿ�A���r���;_��'�?@������R��+~N��<�+~N��R�����?@���'��;_��r���A����ѾQd�F���`   `   )m��[���H澉�;{9���Z��� h�z�4�8m���ؽ�ܮ���
<���󖽏ܮ���ؽ8m�z�4�� h��Z��{9����;H�[���`   `   ���/G���.�־�������y�}��gM��'����Cp��n��]?߽n��Cp������'��gM�y�}��������־�.�/G��`   `   ߦ	�b������t0���ƾ9��v����bp��,Q�)�=�`�3��/���.��/�_�3�)�=��,Q��bp�v���9����ƾt0侼���b��`   `   *��o��o+��"�[�վv�������o��eㅾ���h�������N�����h������eㅾ�o������v��[�վ�"�o+�o��`   `   �������T@���h�T�ɾ���&���;���s���8žо 7Ծо�8ž�s���;��&�����T�ɾ�h�T@������`   `   d�������8�x0�}�ھq�ѾE�־:���t��d����Tz$�����d��t�:��E�־q�Ѿ}�ھx0�8������`   `   k����g�����B���R�쾏���������_<���[�Tt�9}�Tt���[��_<����������R��B������g�����`   `   ���X��9���������������:*�q�U��m�������c��K����c�������m��q�U��:*�������������9��X��`   `   ��|���#��x���,����
��^&�&AW�֩��������!
	�j;�!
	���쿉��֩��&AW��^&���
��,���x���#�|��`   `   8%�Md�2�D�ﾴ���/&��UB��3��찼��|�R�'���F��S���F�R�'��|�찼��3���UB�/&�����D�ﾻ2�Md�`   `   e�վ��վ�a׾!��[����O!��!_��������nG*�LYd��?��ㄕ��?��LYd�nG*�������!_��O!�[���!���a׾��վ`   `   �ʷ� ���[����Ѿ�T���<*��yx�����f��vS���������?����������vS��f�����yx��<*��T����Ѿ�[�� ��`   `   ^������k,������i]����.�;����)ϿJ)!��|s��������N����������|s�J)!��)Ͽ;�����.�i]������k,������`   `   �}�p]��Yt���v��ӷ龻�,�o��uFտf�'�̾����A��*��A�����̾�f�'�uFտo����,�ӷ��v��Yt��p]��`   `   CgK���S��@q�DӘ�2�־2#�J߀�1Ϳ�� �>Us��	�������������	��>Us��� �1ͿJ߀�2#�2�־DӘ��@q���S�`   `   o����'�4*F�A���þ��h��yi�e���b��S��ג�����?������ג��S��b�e���yi��h��þ�A��4*F���'�`   `   ���&;�=��a�Z��C��F���نH�� ����Ǳ)�l>d��E������E��l>d�Ǳ)��뿴 ��نH�F����C��a�Z�=��&;�`   `   ���Cz��k}��R.1��#���*Ӿh~$���z�e��=� ��'�4G�?vS�4G��'�=� �e����z�h~$��*Ӿ�#��R.1�k}��Cz��`   `   b}��z��w��9�� AZ�i���`�(B�����ݻ�"��v�	�G�v�	�"��ݻ�����(B��`�i�� AZ�9��w���z��`   `   �;4�ƅN��/��lO߽��.�$���;˾�h�]�L�Yn������񯼿nWſ񯼿����Yn��]�L��h��;˾$����.�lO߽�/��ƅN�`   `   ���6��">h���������Y��ҟ��?�)��:�A���h�wX��L���wX����h�:�A�)���?��ҟ���Y�������">h�6��`   `   ��Ǽ���>8��N��;�5�9e�����~�������X9��tN�J%V��tN��X9����~������9e��5�;�N���>8����`   `   t�������8�-����ν���*T�Q'�����$��^�>��L��>��^�$�����Q'��*T������ν-����8����`   `   �+��98�m&a�HÔ�Q�ʽ1x
�BJ9�sp�:4��������̾�5޾S侚5޾��̾����:4��sp�BJ9�1x
�Q�ʽHÔ�m&a��98�`   `   !��r���ѝ�yR��_��̼�9�2�ψ^��̆�����H갾�߽��r¾�߽�H갾�����̆�ψ^�9�2�˼�_��yR���ѝ��r��`   `   q��|��.�����t
�$Q�[<��<`�S탾[��-ѧ��޲�?Ķ��޲�-ѧ�[��S탾�<`�[<�$Q��t
�����.��|�`   `   �6=�F];�P7��3�Bx5�	j?��S�Wo�[���L��F��:\�����:\��F��L��Z���Wo��S�	j?�Ax5��3�P7�F];�`   `   Q���:ז������_����w�np�Q�u�0탾<s���Ơ�H���\��Q���\��H����Ơ�<s��0탾Q�u�np���w��_������:ז�`   `   hS��J�t޾7�ž�y��J����$�������1��<a��߲��毽�����毽�߲��<a���1�������$��J����y��7�žt޾J�`   `   �F�a�?��-��3�܀��ξ���秾�ҧ�����_����!���þ�!��_��������ҧ�秾���ξ܀���3��-�a�?�`   `   깝��:���慿��]��0�Y
���޾�b������˳�B��|��5���|��B���˳�����b����޾Y
��0���]��慿�:��`   `   ]���^��AͿ����-#z��Y9��c�L9޾bN��5Ƕ����3����ʹ�3������5Ƕ�bN��L9޾�c��Y9�-#z�����AͿ^��`   `   VsB�]i7�r.�|g���!ev��.�	� ��ϾR8�����W���5Ϯ�W������R8���Ͼ	� ��.�!ev���|g�r.�]i7�`   `   @,������$$f�0�*������'V��j��9޾�Y���ҧ����=Ơ�����ҧ��Y���9޾�j��'V�������0�*�$$f�����`   `   |����J�������i��k��1ȿ���G?(��쾂
���ϝ�[{��/ѐ�[{���ϝ��
����G?(�����1ȿ�k���i�����J��`   `   7�)����<P�������?�����Z9���� ����x��n샾P��n샾�x�� �������Z9������?����<P�����`   `   4�V�C(A�l��ʻ���[����U`��WD�T���jx�������g���]���g����jx��T���WD�U`������[�ʻ��l��C(A�`   `   �ih��Q�����J���#f��	�*���?bF�B���z���Ymp���G��U<���G�Ymp�z���B���?bF�*����	��#f��J������Q�`   `   x�V�*A�i���ͳ�k�[�������WO>�d��V�����R�ʢ(��J�ʢ(���R�V���d��WO>�������k�[��ͳ�i��*A�`   `   ��)�����a��	,��W�?������?-�fZҾ b��Y�3��p
�ab���p
�Y�3� b��fZҾ?-������W�?�	,���a�����`   `   í��K@�������i����ſ�#u�|���䵾ܤa�1y�|Nܽ5KŽ|Nܽ1y�ܤa��䵾|���#u��ſ����i����K@��`   `   ���*����#f���*�9����P�F�~���uۖ�ba9��.��Z��䷔��Z���.�ba9�uۖ�~���P�F���9�쿂�*��#f�*���`   `   ��B�H�7�,E�h��ܬ���k�1_��wþ�}q����ʷ���{�?PX���{��ʷ����}q��wþ1_���k��ܬ�h�,E�H�7�`   `   �����)Tο����2�u��-���ݖ�:�<��潬���28�n8��28������:�<�ݖ����-�2�u�����)Tο��`   `   �������鈿��`�z�,�'7��c)���)g��4�Ҕ��^�Y�N�'��N�^�Y�Ҕ���4��)g�c)��'7��z�,���`�鈿����`   `   J%V��tN��X9����~������9e��5�;�N���>8������Ǽ���>8��N��;�5�9e�����~�������X9��tN�`   `   L��>��^�$�����Q'��*T������ν-����8����t�������8�-����ν���*T�Q'�����$��^�>��`   `   S侚5޾��̾����:4��sp�BJ9�1x
�Q�ʽHÔ�n&a��98��+��98�n&a�HÔ�Q�ʽ1x
�BJ9�sp�:4��������̾�5޾`   `   �r¾�߽�H갾�����̆�ψ^�9�2�̼�_��yR���ѝ��r��"��r���ѝ�yR��_��̼�9�2�ψ^��̆�����H갾�߽�`   `   ?Ķ��޲�-ѧ�[��S탾�<`�[<�$Q��t
�����.��|�q��|��.�����t
�$Q�[<��<`�S탾[��-ѧ��޲�`   `   ���:\��F��L��[���Wo��S�	j?�Bx5��3�P7�F];��6=�F];�P7��3�Bx5�	j?��S�Wo�[���L��F��:\��`   `   Q���\��H����Ơ�<s��0탾Q�u�np���w��_������:ז�Q���:ז������_����w�np�Q�u�0탾<s���Ơ�H���\��`   `   ����毽�߲��<a���1�������$��J����y��7�žt޾J�hS��J�t޾7�ž�y��J����$�������1��<a��߲��毽�`   `   �þ�!��_��������ҧ�秾���ξ܀���3��-�a�?��F�a�?��-��3�܀��ξ���秾�ҧ�����_����!��`   `   5���|��B���˳�����b����޾Y
��0���]��慿�:��깝��:���慿��]��0�Y
���޾�b������˳�B��|��`   `   �ʹ�3������5Ƕ�bN��L9޾�c��Y9�-#z�����AͿ^��]���^��AͿ����-#z��Y9��c�L9޾bN��5Ƕ����3���`   `   5Ϯ�W������R8���Ͼ	� ��.�!ev���|g�r.�]i7�VsB�]i7�r.�|g���!ev��.�	� ��ϾR8�����W���`   `   =Ơ�����ҧ��Y���9޾�j��'V�������0�*�$$f�����@,������$$f�0�*������'V��j��9޾�Y���ҧ����`   `   /ѐ�[{���ϝ��
����G?(�����1ȿ�k���i�����J��|����J�������i��k��1ȿ���G?(��쾂
���ϝ�[{��`   `   P��n샾�x�� �������Z9������?����<P�����7�)����<P�������?�����Z9���� ����x��n샾`   `   ��]���g����jx��T���WD�U`������[�ʻ��l��C(A�4�V�C(A�l��ʻ���[����U`��WD�T���jx�������g�`   `   �U<���G�Ymp�z���B���?bF�*����	��#f��J������Q��ih��Q�����J���#f��	�)���?bF�A���z���Ymp���G�`   `   �J�ʢ(���R�V���d��WO>�������k�[��ͳ�i��*A�x�V�*A�i���ͳ�j�[�������WO>�d��V�����R�ʢ(�`   `   ab���p
�Y�3� b��fZҾ?-������W�?�	,���a�������)�����a��	,��W�?������?-�fZҾ b��Y�3��p
�`   `   5KŽ|Nܽ1y�ܤa��䵾|���#u��ſ����i����K@��í��K@�������i����ſ�#u�|���䵾ܤa�1y�|Nܽ`   `   ䷔��Z���.�ba9�uۖ�~���P�F���9�쿂�*��#f�*������*����#f���*�9����P�F�~���uۖ�ba9��.��Z��`   `   ?PX���{��ʷ����}q��wþ1_���k��ܬ�h�,E�H�7���B�H�7�,E�h��ܬ���k�1_��wþ�}q����ʷ���{�`   `   n8��28������:�<�ݖ����-�2�u�����)Tο�����)Tο����2�u��-���ݖ�:�<��潬���28�`   `   '��N�^�Y�Ҕ���4��)g�c)��'7��z�,���`�鈿�����������鈿��`�z�,�'7��c)���)g��4�Ҕ��^�Y�N�`   `   N��~ڼ�d,��u��5���C5�aۆ������~��%��&G�@_�,h�@_��&G��%��~�����aۆ��C5�5���u���d,�~ڼ`   `   %Ӽ]����&�:�z�I����<�
}H������=���_�����������������_ྏ=������
}H��<�H���:�z���&�]��`   `   m�"��c,���K�+R������+l�e����Q�Q���]���B����ɾ��Ͼ��ɾB��]���Q�����Q�e��+l�����+R����K��c,�`   `   Zx������$㓽����g��ٓ彲=�(0�&�U��n{�
���!ܘ�����!ܘ�
����n{�&�U�(0��=�ؓ彗g�����$㓽����`   `   �x�y�����e罷e� 8���i���%���?�TZ��q��؀�廙��؀��q�TZ���?���%��i� 8���e�e����y��`   `   :FJ��IF�W�;���.��b#�!��� ���+�o�<�&P���a�
hn���r�
hn���a�&P�o�<���+��� �!��b#���.�W�;��IF�`   `   ݲ����������ֆ��l��Q���B���?�NgF��R�0
`�J�i��m�J�i�0
`��R�NgF���?���B��Q��l��ֆ��������`   `   f�
��=��)vѾ�K��)l�� �v���_���X�$7\��Ed�L�k�Zn�L�k��Ed�$7\���X���_� �v�)l���K��)vѾ��=�`   `   omb�M�Y��(B��P"�y}�\vʾ%���zK��;�q�i�y�i���m��]o���m�y�i�i�;�q�zK��%���\vʾy}��P"��(B�M�Y�`   `   �����^��W���R�y��?�$����Ӿ1��v���"�w���n��xm���m��xm���n�!�w�v���1����Ӿ$���?�R�y�W����^��`   `   �]�����M���1`���'G������ɾ�ț�������q�@�i�Ch�@�i���q������ț���ɾ����'G�1`�����M����`   `   ��p���a��;��S��~ɿۣ��&V6������ر�g싾��r�c&c��_�c&c���r�g싾�ر�����&V6�ۣ���~ɿ�S��;���a�`   `   5���Ŵ�����UP�vc�����>h�<��-�ɾ�(����q�{Y��R�{Y���q��(��-�ɾ<��>h�����vc�UP����Ŵ��`   `   Ns$�1t�[�����;�Ii�wh����/�X�h���F�n�ψM��D�ψM�E�n�h���X���/�wh��Ii迗�;��[��1t�`   `   ��s��g[��1 �����W(l�Wc������'G�$��g��� �h���?���3���?� �h�g���$���'G�����Wc�W(l������1 ��g[�`   `   )̚��C��x�J�N����n���`�,ѷ��W�=� ������_���/�""���/���_����=� ��W�,ѷ��`��n��N���x�J��C��`   `   �����Ö��g[������H-%����!\�/}�;d����Q�8p�0[�8p���Q�;d��/}��!\���H-%�������g[��Ö�`   `   �˚�sE��|�J����G�����������T�����e-���)?�3�:���3��)?�e-�������T��������G������|�J�sE��`   `   (�s��g[�D �����l�>���ڥ��)B���Ն� m(��M�J�Ͻ�M� m(�Ն����)B��ڥ�>���l����D ��g[�`   `   l^$�@i�c!���Г�<�����ӌ���'�l�ž7wi����-ý�ا�-ý���7wi�l�ž��'��ӌ����<��Г�c!��@i�`   `   ����e�������P�s��_p��(pb�"�	�����A����C7���;��C7������A����"�	�(pb�_p��s���P����e���`   `   �p��a��;��j��^ɿ���!�-��Wؾ����\�������i��A���i������\�����Wؾ!�-�����^ɿ�j��;��a�`   `   [��c�f&�k��r����+B��� �����FI�g|�����HR,��`�HR,�����g|FI������ ��+B�r���k��f&�c�`   `   �������8f��Ǯz�_>����8���ݳs��<������S�� �J�ͼ� ���S�����<�ݳs�8������_>�Ǯz�8f������`   `   ,h�@_��&G��%��~�����aۆ��C5�5���u���d,�~ڼN��~ڼ�d,��u��5���C5�aۆ������~��%��&G�@_�`   `   ����������_ྏ=������
}H��<�I���:�z���&�^��%Ӽ^����&�:�z�I����<�
}H������=���_�������`   `   ��Ͼ��ɾB��]���Q�����Q�e��+l�����+R����K��c,�m�"��c,���K�+R������+l�e����Q�Q���]���B����ɾ`   `   ����!ܘ�
����n{�&�U�(0��=�ٓ彗g�����$㓽����Zx������$㓽����g��ٓ彲=�(0�&�U��n{�
���!ܘ�`   `   廙��؀��q�TZ���?���%��i� 8���e�e����y���x�y�����e罷e� 8���i���%���?�TZ��q��؀�`   `   ��r�
hn���a�&P�o�<���+��� �!��b#���.�W�;��IF�:FJ��IF�W�;���.��b#�!��� ���+�o�<�&P���a�
hn�`   `   �m�J�i�0
`��R�NgF���?���B��Q��l��ֆ��������ݲ����������ֆ��l��Q���B���?�NgF��R�0
`�J�i�`   `   Zn�L�k��Ed�$7\���X���_� �v�)l���K��)vѾ��=�f�
��=��)vѾ�K��)l�� �v���_���X�$7\��Ed�L�k�`   `   �]o���m�y�i�i�;�q�zK��%���\vʾy}��P"��(B�M�Y�omb�M�Y��(B��P"�y}�\vʾ%���zK��;�q�i�y�i���m�`   `   ��m��xm���n�"�w�v���1����Ӿ$���?�R�y�W����^�������^��W���R�y��?�$����Ӿ1��v���!�w���n��xm�`   `   Ch�@�i���q������ț���ɾ����'G�1`�����M�����]�����M���1`���'G������ɾ�ț�������q�@�i�`   `   �_�c&c���r�g싾�ر�����&V6�ۣ���~ɿ�S��;���a���p���a��;��S��~ɿۣ��&V6������ر�g싾��r�c&c�`   `   �R�{Y���q��(��-�ɾ<��>h�����vc�UP����Ŵ��5���Ŵ�����UP�vc�����>h�<��-�ɾ�(����q�{Y�`   `   �D�ψM�F�n�h���X���/�wh��Ii迗�;��[��1t�Ns$�1t�[�����;�Ii�wh����/�X�h���E�n�ψM�`   `   ��3���?� �h�g���$���'G�����Wc�W(l������1 ��g[���s��g[��1 �����W(l�Wc������'G�$��g��� �h���?�`   `   ""���/���_����=� ��W�,ѷ��`��n��N���x�J��C��)̚��C��w�J�N����n���`�,ѷ��W�=� ������_���/�`   `   0[�8p���Q�;d��/}��!\���H-%�������g[��Ö������Ö��g[������H-%����!\�/}�;d����Q�8p�`   `   :���3��)?�e-�������T��������G������|�J�sE���˚�sE��|�J����G�����������T�����e-���)?�3�`   `   J�Ͻ�M� m(�Ն����)B��ڥ�>���l����D ��g[�(�s��g[�D �����l�>���ڥ��)B���Ն� m(��M�`   `   �ا�-ý���7wi�l�ž��'��ӌ����<��Г�c!��@i�l^$�@i�c!���Г�<�����ӌ���'�l�ž7wi����-ý`   `   �;��C7������A����"�	�(pb�_p��s���P����e�������e�������P�s��_p��(pb�"�	�����A����C7��`   `   �A���i������\�����Wؾ!�-�����^ɿ�j��;��a��p��a��;��j��^ɿ���!�-��Wؾ����\�������i�`   `   �`�HR,�����g|FI������ ��+B�r���k��f&�c�[��c�f&�k��r����+B��� �����FI�g|�����HR,�`   `   J�ͼ� ���S�����<�ݳs�8������_>�Ǯz�8f�������������8f��Ǯz�_>����8���ݳs��<������S�� �`   `   P����%ͼ�a$�������㽥'3�╆������k�F)�K�L�Xf��no�Xf�K�L�F)��k�����╆��'3���㽓����a$��%ͼ`   `   �ƼW�Z��$�g�?K��4���>>�����ٵ��B`۾�����?9������B`۾ٵ�������>>�4��?K��$�g�Z��W�`   `   8���c$�<�<��bj��@��ݴн.��;��*o��4��߰��w����п�w���߰���4���*o��;�.�ݴн�@���bj�<�<��c$�`   `   \d��E։� D��甓�񅣽�q�������/��+O��Lk���~�-Ƃ���~��Lk��+O��/����齇q��񅣽甓� D��E։�`   `   j��W�����!ؽ,�н܃ҽ^�ཛྷ���R����!���2��>�$C��>���2���!�R������^��܃ҽ,�н�!ؽ��W��`   `   �_P��K�a�<�)����^���������������������!��������������������^���)�a�<��K�`   `   ԯ��V��OT��l���0Ma�x;�������s��G	�Xd�h���h�Xd��G	��s������x;�0Ma�l���OT���V��`   `   �
�+���1��"�վ�=��p����T��c.�{��b$�o��Li�G��Li�o��b$�{���c.���T�p���=��"�վ�1��+��`   `   p�pf�_AL���(�`j�%ž|5��Y^���2����Ch�`��J�_��Ch������2�Y^�|5��%ž`j���(�_AL�pf�`   `   bĿ8]��Y������F�N���ɾG�����V��g-�ܐ����6����ܐ��g-���V�G�����ɾN�F�����Y��8]��`   `   �� ���m���ʿ񅓿ԉL���	�����聾�C�q!�Cd���Cd�q!��C�聾������	�ԉL�񅓿�ʿm����`   `   jτ�0x���L�v���qֿ~�����8�q�u���c�[��*�.��i��.���*�c�[�u���q��8�~����qֿv����L�0x�`   `   ����Y��<ǡ��d�H(������oo�������ZTv�r�2�����<	����r�2�ZTv��������oo�����H(��d�<ǡ��Y��`   `   @�C�,�'_�������:L�N���㔿��1�|<׾�ч�5`:�N{� w�N{�5`:��ч�|<׾��1��㔿N���:L�����'_��C�,�`   `   �ߎ�o~����:�ǭ�����*(�
ů���L�^��/���@?�o���8 �o���@?��/��^����L�
ů�*(����ǭ����:�o~��`   `   �:��?��lHm�\������Kp+�6.ÿVB_�9� ��Z����?�)]	�rt�)]	���?��Z��9� �VB_�6.ÿKp+�����\��lHm�?��`   `   
���{��o~����)ǡ��:3��ʿ�f��h�����:��M��UབM���:����h��f��ʿ�:3�)ǡ���o~��{��`   `   �9��1
��(Ym���Q��A�+�T�ÿ'X_�6���챒���/��^�(�ɽ�^콄�/�챒�6���'X_�T�ÿA�+�Q����(Ym�1
��`   `   �ڎ�t~���;����*�����&ְ�BL�1\��c���нu����нc���1\�BL�&ְ���*�������;�t~��`   `   ��?���,����A"��fVM��M��/ٕ��|0���̾�k�̏	�ס���Œ�ס��̏	��k���̾�|0�/ٕ��M��fVM�A"�������,�`   `   �������]ǡ�E�d�/��¿�!p����|W��i�D�N�㽭����$j�����N��i�D�|W������!p��¿/�E�d�]ǡ����`   `   �G��"Yw���L�Y����׿�u��!i7�r��l��2�@����\�E�1���\�@��2�l��r��!i7��u����׿Y����L�"Yw�`   `   D��%(��?�ψʿ�蓿jDL����[���O�����s���I$�%���I$��s�����O�[�����jDL��蓿ψʿ�?�%(�`   `   [�¿��������Db���dF��s�;鿾Ѫx�{��̺����N����:������N�̺��{��Ѫx�;鿾�s��dF�Db����������`   `   �no�Xf�K�L�F)��k�����╆��'3���㽓����a$��%ͼP����%ͼ�a$�������㽥'3�╆������k�F)�K�L�Xf�`   `   ?9������B`۾ٵ�������>>�4��?K��$�g�Z��W��ƼW�Z��$�g�?K��4���>>�����ٵ��B`۾�����`   `   �п�x���߰���4���*o��;�.�ݴн�@���bj�<�<��c$�8���c$�<�<��bj��@��ݴн.��;��*o��4��߰��x���`   `   -Ƃ���~��Lk��+O��/����齇q��񅣽甓� D��E։�\d��E։� D��甓�񅣽�q�������/��+O��Lk���~�`   `   $C��>���2���!�R������^��܃ҽ,�н�!ؽ��W��j��W�����!ؽ,�н܃ҽ^�ཛྷ���R����!���2��>�`   `   ��!��������������������^���)�a�<��K��_P��K�a�<�)����^�������������������`   `   ��h�Xd��G	��s������x;�0Ma�l���OT���V��ԯ��V��OT��l���0Ma�x;�������s��G	�Xd�h�`   `   G��Li�o��b$�{���c.���T�p���=��"�վ�1��+���
�+���1��"�վ�=��p����T��c.�{��b$�o��Li�`   `   J�`��Ch������2�Y^�|5��%ž`j���(�_AL�pf�p�pf�_AL���(�`j�%ž|5��Y^���2����Ch�`��`   `   6����ܐ��g-���V�G�����ɾN�F�����Y��8]��bĿ8]��Y������F�N���ɾG�����V��g-�ܐ����`   `   ��Cd�q!��C�聾������	�ԉL�񅓿�ʿm������ ���m���ʿ񅓿ԉL���	�����聾�C�q!�Cd�`   `   i��.���*�c�[�u���q��8�~����qֿv����L�0x�jτ�0x���L�v���qֿ~�����8�q�u���c�[��*�.��`   `   �<	����r�2�ZTv��������oo�����H(��d�<ǡ��Y������Y��<ǡ��d�H(������oo�������ZTv�r�2����`   `    w�N{�5`:��ч�|<׾��1��㔿N���:L�����'_��C�,�@�C�,�'_�������:L�N���㔿��1�|<׾�ч�5`:�N{�`   `   �8 �o���@?��/��^����L�
ů�*(����ǭ����:�o~���ߎ�o~����:�ǭ�����*(�
ů���L�^��/���@?�o��`   `   qt�)]	���?��Z��9� �VB_�6.ÿKp+�����]��lHm�?���:��?��lHm�\������Kp+�6.ÿVB_�9� ��Z����?�)]	�`   `   �UབM���:����h��f��ʿ�:3�)ǡ���o~��{��
���{��o~����)ǡ��:3��ʿ�f��h�����:��M�`   `   (�ɽ�^콄�/�챒�6���'X_�T�ÿA�+�Q����(Ym�1
���9��1
��'Ym���Q��A�+�T�ÿ'X_�6���챒���/��^�`   `   u����нb���1\�BL�&ְ���*�������;�t~���ڎ�t~���;����*�����&ְ�BL�1\��b���н`   `   �Œ�ס��̏	��k���̾�|0�/ٕ��M��fVM�A"�������,���?���,����A"��fVM��M��/ٕ��|0���̾�k�̏	�ס��`   `   �$j�����N��i�D�|W������!p��¿/�E�d�]ǡ�����������]ǡ�E�d�/��¿�!p����|W��i�D�N�㽭���`   `   E�1���\�@��2�l��r��!i7��u����׿Y����L�"Yw��G��"Yw���L�Y����׿�u��!i7�r��l��2�@����\�`   `   %���I$��s�����O�[�����jDL��蓿ψʿ�?�%(�D��%(��?�ψʿ�蓿jDL����[���O�����s���I$�`   `   :������N�̺��{��Ѫx�;鿾�s��dF�Db����������[�¿��������Db���dF��s�;鿾Ѫx�{��̺����N����`   `   3����㾼�F�T����ؽP+�G〾�2�������#��#E���]�x�f���]��#E��#������2��G〾P+���ؽT���F��㾼`   `   N����Ѽ���*�T�>��c.󽁴0��v�Xq�ξW7��MA�?4�MA�W7��q�ξX�v���0�c.�>��+�T�����Ѽ`   `   U��bJ�mJ-���R����Z෽af��X0&�� V�������.���L6��.���������� V�X0&�af��Z෽�����R�mJ-�bJ�`   `   ����������� ��~!�����H���+��H�-�,�oE��wV�В\��wV�oE�-�,�H�+��H������~!�� ����������`   `   뽛��{ؽ"&ǽ�ڷ�#����ⲽ�
��8-ؽa�����$�y�$����a��8-ؽ�
���ⲽ#����ڷ�"&ǽ{ؽ���`   `   D�K��E�'�5�PB�-���<潗�ɽo����E���U��8�˽�?Խۉ׽�?Խ8�˽�U���E��o�����ɽ�<�-��PB�'�5��E�`   `   �}��{¦������ހ�@�Q��,&����-ؽ6��!��N[��b8���b8��N[��!��6���-ؽ���,&�@�Q��ހ�����{¦�`   `   �L��
�\+����ξ����x��S8��v
���ٽ�D��%�������K������%����D����ٽ�v
��S8��x������ξ\+���
�`   `   T>k��a�W�G�x�#�����5Y��)���5�9�����pн�6��|���A��|����6���pн���5�9�)���5Y������x�#�W�G��a�`   `   �ֿ�����z��!��.A@�I��R����{�P�+�����ܿ�����ǝ������ܿ����P�+���{�R��I��.A@�!���z�����`   `   EQ�f��Þ���9ſmR���#E�5\�A����[��v�s�ֽ�+���o���+��s�ֽ�v��[�A���5\��#E�mR���9ſÞ��f��`   `   Wc���%p�n�F��/��qп�7��]�0�h�ܾ���� $0��Z�����F������Z� $0�����h�ܾ]�0��7���qп�/�n�F��%p�`   `   �$��|���ʛ���\����ݺ���f����t����O�E��Pƽ���PƽE���O�t��������f�ݺ������\�ʛ�|���`   `   M�6��$�u���a�����E�#%�5���**�C�Ǿ�im�P7�'�н�}��'�нP7��im�C�Ǿ�**��5��#%��E�a���u����$�`   `   :͇�^8t���1������H{��������k"E����c�����s ؽjt��s ؽ��c������k"E���������H{�������1�^8t�`   `   <G��s ��za� ?�m4���f&��ѽ�:@X����A��?�%�zSڽ���zSڽ?�%�A�����:@X��ѽ��f&�m4�� ?�za�s ��`   `   #����ȧ�q8t�@��5ʛ�E�-��9ſ��_�{���� ��!&��ֽ����ֽ!&�� ��{�����_��9ſE�-�5ʛ�@��q8t��ȧ�`   `   �F�����C�a��`������'�L���y�Y�����k��]��,nʽ���,nʽ]��k������y�Y�L����'������`�C�a����`   `   ȇ��8t�	�1�%��w|�������G���㾼؀��*�+����-��+����*��؀�����G������w|�%��	�1��8t�`   `   �z6�cq$�p���;���l7G�u��V�����,���ǾaBc��E��/���耽�/���E�aBc���Ǿ��,�V���u��l7G�;���p���cq$�`   `   ����1U��xʛ�	�]�{��L���}Ak�c���¦��>�#bؽTD���@R�TD��#bؽ�>��¦�c��}Ak�L���{��	�]�xʛ�1U��`   `   ��X'o�WF����,;ҿ&N����3��G޾������\�����M�]p"���M�\����������G޾��3�&N��,;ҿ���WF�X'o�`   `   �����UL���:ſ?N����G�u���Ʀ�D_J�q�$都s*�K��s*�$都q�D_J��Ʀ�u����G�?N���:ſUL����`   `   g�����������]�Z�@���	�7����q���y,��hvE�	�弃���	��hvE�y,�����q�7�����	�Z�@��]���������`   `   x�f���]��#E��#������2��G〾P+���ؽT���F��㾼3����㾼�F�T����ؽP+�G〾�2�������#��#E���]�`   `   ?4�MA�W7��q�ξX�v���0�c.�>��+�T�����ѼO����Ѽ���+�T�>��c.󽁴0��v�Xq�ξW7��MA�`   `   L6��.���������� V�X0&�af��Z෽�����R�nJ-�bJ�U��bJ�nJ-���R����Z෽af��X0&�� V�������.���`   `   В\��wV�oE�-�,�H�+��H������~!�� ��������������������� ��~!�����H���+��H�-�,�oE��wV�`   `   y�$����a��8-ؽ�
���ⲽ#����ڷ�"&ǽ{ؽ���뽛��{ؽ"&ǽ�ڷ�#����ⲽ�
��8-ؽa�����$�`   `   ۉ׽�?Խ8�˽�U���E��o�����ɽ�<�-��QB�'�5��E�D�K��E�'�5�PB�-���<潗�ɽo����E���U��8�˽�?Խ`   `   �b8��N[��!��6���-ؽ���,&�@�Q��ހ�����{¦��}��{¦������ހ�@�Q��,&����-ؽ6��!��N[��b8��`   `   K������%����D����ٽ�v
��S8��x������ξ\+���
��L��
�\+����ξ����x��S8��v
���ٽ�D��%�������`   `   A��|����6���pн���5�9�)���5Y������x�#�W�G��a�T>k��a�W�G�x�#�����5Y��)���5�9�����pн�6��|���`   `   ǝ������ܿ����P�+���{�R��I��.A@�!���z������ֿ�����z��!��.A@�I��R����{�P�+�����ܿ�����`   `   �o���+��s�ֽ�v��[�A���5\��#E�mR���9ſÞ��f��EQ�f��Þ���9ſmR���#E�5\�A����[��v�s�ֽ�+��`   `   �F������Z� $0�����h�ܾ]�0��7���qп�/�n�F��%p�Wc���%p�n�F��/��qп�7��]�0�h�ܾ���� $0��Z����`   `   ���PƽE���O�t��������f�ݺ������\�ʛ�|����$��|���ʛ���\����ݺ���f����t����O�E��Pƽ`   `   �}��'�нP7��im�C�Ǿ�**��5��#%��E�a���u����$�M�6��$�u���a�����E�#%�5���**�C�Ǿ�im�P7�'�н`   `   jt��s ؽ��c������k"E���������H{�������1�^8t�:͇�^8t���1������H{��������k"E����c�����s ؽ`   `   ���zSڽ?�%�A�����:@X��ѽ��f&�m4�� ?�za�s ��<G��s ��za� ?�m4���f&��ѽ�:@X����A��?�%�zSڽ`   `   ����ֽ!&�� ��{�����_��9ſE�-�5ʛ�@��q8t��ȧ�#����ȧ�q8t�@��5ʛ�E�-��9ſ��_�{���� ��!&��ֽ`   `   ���,nʽ]��k������y�Y�L����'������`�C�a�����F�����C�a��`������'�L���y�Y�����k��]��,nʽ`   `   �-��+����*��؀�����G������w|�%��	�1��8t�ȇ��8t�	�1�%��w|�������G���㾼؀��*�+���`   `   �耽�/���E�aBc���Ǿ��,�V���u��l7G�;���p���cq$��z6�cq$�p���;���l7G�u��V�����,���ǾaBc��E��/��`   `   �@R�TD��#bؽ�>��¦�c��}Ak�L���{��	�]�xʛ�1U������1U��xʛ�	�]�{��L���}Ak�c���¦��>�#bؽTD��`   `   ]p"���M�\����������G޾��3�&N��,;ҿ���WF�X'o���X'o�WF����,;ҿ&N����3��G޾������\�����M�`   `   K��s*�$都q�D_J��Ʀ�u����G�?N���:ſUL���������UL���:ſ?N����G�u���Ʀ�D_J�q�$都s*�`   `   ����	��hvE�y,�����q�7�����	�Z�@��]���������g�����������]�Z�@���	�7����q���y,��hvE�	��`   `   :v������&
���l�suĽ�U���i�Q����W侲����0�F�F�ְN�F�F���0�����W�Q�����i��U�suĽ��l�&
�����`   `   �[�������	��6s<��叽�{ؽɥ�+3\�倒�����C�ھ7�,���7�C�ھ����倒�+3\�ɥ��{ؽ�叽6s<��	������`   `   ��3+
��-��7�'�k��h��Y(׽r����9�?Me������h���>���h������?Me���9�r��Y(׽�h��'�k��7��-�3+
�`   `   �lq��,o��j��i��]r�Ć�g��oý���q��1�#��2�aM7��2�1�#�q�����oýg��Ć��]r��i��j��,o�`   `   �Xؽ��ҽ�mĽ
���b������#�� ͔�����N跽�˽?�ٽZ2߽?�ٽ�˽N跽���� ͔��#������b��
���mĽ��ҽ`   `   ��;��6��&�~�c(�f/½�������B9��k��G\��6틽�΍�6틽G\��k��B9���������f/½c(�~��&��6�`   `   у�����&����i�Z;����7(ؽ�����Q���_��M��%G�_�E��%G��M��_��Q������7(ؽ���Z;���i��&����`   `   [������l���-e���[��u�D۽[e���[g�}�:�UC%���UC%�}�:��[g�[e��D۽�u��[�-e�����l����`   `   6�T��!L���4���1S������Ke������˽�щ��G��} �����} ��G��щ���˽����Ke�����1S�����4��!L�`   `   `#���w��J㎿�mf�=5-��c��͉��J$W��������i���-�u
���-��i�������J$W�͉���c��=5-��mf�J㎿�w��`   `   +�����V�޿�d��rM����0�����g����5�(߽BC��uG�|�-�uG�BC��(߽��5��g����辫�0�rM���d��V�޿���`   `   n|Z��DM���+�l���Ӹ�(.w��7��þ4�k��p��"���f��E��f��"���p�4�k��þ�7�(.w��Ӹ�l����+��DM�`   `   ����XM��~o��q�=�� ����N�����d��;�+��w˽p΄���^�p΄��w˽;�+��d������N���� �q�=�~o��XM��`   `   p��g �ֶ��[y����*�ӸԿ�Ѐ�!s�7ڰ�^�J�U 뽺���˜w�����U �^�J�7ڰ�!s��Ѐ�ӸԿ��*�[y��ֶ��g �`   `   1KQ�F<�(/
��F����U�� ����T�0��ʾ�:e����ģ�����ģ����:e��ʾT�0����� ���U��F��(/
�F<�`   `   ���K o���-����h�w���!Ԩ�eB�~�ܾ��w��>������������>���w�~�ܾeB�!Ԩ���h�w������-�K o�`   `   ��Ym��5F<������o���f�9e���fI�iN侌��Z���z䍽�Z�����iN侲fI�9e���f��o������5F<�Ym��`   `   ��fo��.�����'Qx����.��R�D���߾�z�\��v����,��v���\���z���߾R�D��.����'Qx������.�fo�`   `   }AQ�OF<�]H
�����7W����Yz����4���Ͼ<�i�%�@0����|�@0��%�<�i���Ͼ��4�Yz�����7W�����]H
�OF<�`   `   W��@X ��������H,���׿�˃�+*��ܶ��}O�n���Y��oj]��Y��n���}O��ܶ�+*��˃���׿�H,�������@X �`   `   ;G��� ��p��=K>�E��u0���T���q��#/��RĽ��h�r87���h��RĽ#/�q�����T�u0��E��=K>�p��� ��`   `   eAY�"GL�
d+���ֺ��{|��q#�ٰ˾OXt����(]���7�����7�(]�����OXt�ٰ˾�q#��{|�ֺ���
d+�"GL�`   `   W�}� �x�ݿ�f������4�>������n:�fUؽK�p�	
���Ӽ	
�K�p�fUؽ�n:����>���4�����f��x�ݿ}� �`   `   
駿���=���Ae�P;.�)���oh���c]����g��X/3���̼xz����̼X/3�g������c]�oh��)���P;.��Ae�=�����`   `   ְN�F�F���0�����W�Q�����i��U�suĽ��l�&
�����;v������&
���l�suĽ�U���i�Q����W侲����0�F�F�`   `   ,���7�C�ھ����倒�+3\�ɥ��{ؽ�叽6s<��	�������[�������	��6s<��叽�{ؽɥ�+3\�倒�����C�ھ7�`   `   �>���h������?Me���9�r��Y(׽�h��'�k��7��-�4+
���3+
��-��7�'�k��h��Y(׽r����9�?Me������h��`   `   aM7��2�1�#�q�����oýg��Ć��]r��i��j��,o��lq��,o��j��i��]r�Ć�g��oý���q��1�#��2�`   `   Z2߽?�ٽ�˽N跽���� ͔��#������b��
���mĽ��ҽ�Xؽ��ҽ�mĽ
���b������#�� ͔�����N跽�˽?�ٽ`   `   �΍�6틽G\��k��B9���������f/½d(�~��&��6���;��6��&�~�c(�f/½�������B9��k��G\��6틽`   `   _�E��%G��M��_��Q������7(ؽ���Z;���i��&����у�����&����i�Z;����7(ؽ�����Q���_��M��%G�`   `   ��UC%�}�:��[g�[e��D۽�u��[�-e�����l����[������l���-e���[��u�D۽[e���[g�}�:�UC%�`   `   ����} ��G��щ���˽����Ke�����1S�����4��!L�6�T��!L���4���1S������Ke������˽�щ��G��} �`   `   u
���-��i�������J$W�͉���c��=5-��mf�J㎿�w��`#���w��J㎿�mf�=5-��c��͉��J$W��������i���-�`   `   |�-�uG�BC��(߽��5��g����辫�0�rM���d��V�޿���+�����V�޿�d��rM����0�����g����5�(߽BC��uG�`   `   �E��f��"���p�4�k��þ�7�(.w��Ӹ�l����+��DM�n|Z��DM���+�l���Ӹ�(.w��7��þ4�k��p��"���f�`   `   ��^�p΄��w˽;�+��d������N���� �q�=�~o��XM������XM��~o��q�=�� ����N�����d��;�+��w˽p΄�`   `   ˜w�����U �^�J�7ڰ�!s��Ѐ�ӸԿ��*�[y��ֶ��g �p��g �ֶ��[y����*�ӸԿ�Ѐ�!s�7ڰ�^�J�U 뽺���`   `   ����ģ����:e��ʾT�0����� ���U��F��(/
�F<�1KQ�F<�(/
��F����U�� ����T�0��ʾ�:e����ģ�`   `   ��������>���w�~�ܾeB�!Ԩ���h�w������-�K o����K o���-����h�w���!Ԩ�eB�~�ܾ��w��>����`   `   z䍽�Y�����iN侲fI�9e���f��o������5F<�Ym����Ym��5F<������o���f�9e���fI�iN侌��Y���`   `   �,��v���\���z���߾R�D��.����'Qx������.�fo���fo��.�����'Qx����.��R�D���߾�z�\��v���`   `   ��|�@0��%�<�i���Ͼ��4�Yz�����7W�����]H
�OF<�}AQ�OF<�]H
�����7W����Yz����4���Ͼ<�i�%�@0��`   `   oj]��Y��n���}O��ܶ�+*��˃���׿�H,�������@X �W��@X ��������H,���׿�˃�+*��ܶ��}O�n���Y��`   `   r87���h��RĽ#/�q�����T�u0��E��=K>�p��� ��;G��� ��p��=K>�E��u0���T���q��#/��RĽ��h�`   `   ����7�']�����OXt�ٰ˾�q#��{|�ֺ���
d+�"GL�eAY�"GL�
d+���ֺ��{|��q#�ٰ˾OXt����(]���7�`   `   ��Ӽ	
�K�p�fUؽ�n:����>���4�����f��x�ݿ}� �W�}� �x�ݿ�f������4�>������n:�fUؽK�p�	
�`   `   xz����̼X/3�g������c]�oh��)���P;.��Ae�=�����
駿���=���Ae�P;.�)���oh���c]����g��X/3���̼`   `   ��Q��䆼8_���H�����Z���G�+�������������q%���+��q%����������+�����G�Z�������H�9_��䆼`   `   ^u������Q�μ�����q�ֶ��`��-:� 7w��R��{����˾��Ҿ�˾{����R�� 7w��-:��`�ֶ���q����Q�μ����`   `   X�޼�h��������A�y�������/�� �{J>��]^���t�\�|���t��]^�{J>�� ��/���y����A�������h�`   `   �;N���K�ٟE�w]A�E�w?X���}��͚��뽽Z��p�����~�����p��Z���뽽�͚���}�w?X�E�w]A�ٟE���K�`   `   պ�~�����g5��Ms���th�YJ[��{_�(�r��}�����F󠽣���F󠽴���}��(�r��{_�YJ[��th�Ms��g5����~���`   `   cm"�^6�����{���\ǽ�Z�x�b�K�e�3��+�T�,�F�0�,�2�F�0�T�,��+�e�3�b�K�Z�x���\ǽ�{�����^6�`   `   �F��.����m���G��}��&����+�r���-�E��`�ڼ��ż�'����ż`�ڼE����-�+�r�����&}���G��m�.���`   `   p�޾r־�����(���z��7��6��8��W��L������n��zWe��n�������L��W�8��6���7��z��(������r־`   `   �(2��*+�	��������ߍ���F>��k������.�C�żul�I\;�ul�C�ż�.�����k���F>�ߍ���������	��*+�`   `   �`��I[���,l���?�:3�zeξ����40�Z�ӽ��p�[���*��ƘZ��*��[����p�Z�ӽ40�����zeξ:3���?��,l�I[��`   `   Cڿ��Ͽ���n`��{dT�����þܤt����$礽�2��ż����ż�2�$礽���ܤt��þ���{dT�n`�������Ͽ`   `   �m'�aA��B�пF���W�L��>��j���A���ٽ�Rl����fʼ���Rl���ٽ�A��j���>�W�L�F���B�п�aA�`   `   ��|�'�l���C����jͿI·���+�2Ѿ��t�}|	����+�����+���}|	���t�2Ѿ��+�I·��jͿ����C�'�l�`   `   ���O���פ��pF����@ث�e�T����䓾̬%�C��w�P��"�w�P�C��̬%�䓾���e�T�@ث����pF�פ��O���`   `   uW�%���n��*C|�!$�kͿ>�y�t���<���5>�
�нSDr�/�<�SDr�
�н�5>��<��t��>�y�kͿ!$�*C|��n��%��`   `   �R&����������:�����$��uV"��#����O�o佪^��J�P��^��o���O��#��uV"��$�������:��������`   `   F�3��"�s%��������C��h�Ka���J(�1��r�W����t����Z��t����r�W�1���J(�Ka���h���C�����s%���"�`   `   �Q&��
��������-�;�H翄s��K�$�����U���뽠n��\WY��n�����U�����K�$��s��H�-�;���������
�`   `   pO��%��陷�S�|�9%���Ͽ��~��
�5ٰ�M�G���ݽ@���HL�@����ݽM�G�5ٰ��
���~���Ͽ9%�S�|�陷��%��`   `   �Q��W����ŉ�T=G�S���Ӯ���Z����+s���$2��ƽ��g��5���g��ƽ�$2�,s�������Z��Ӯ�S��T=G��ŉ�W���`   `   8D|��l�^�C������Ͽ�ڊ�T-2�B�ܾ������J֧��B�2���B�J֧�������B�ܾT-2��ڊ���Ͽ���^�C��l�`   `   3V&��_�v)�Usѿ�n����Q�p
�@K���R�|N󽷹��H�����H������|N��R�@K��p
���Q��n��Usѿv)��_�`   `    z׿=lͿF����b��@�V���>�̾f���}!��Ѻ�qtM�Q%�ޫ�Q%�qtM��Ѻ�}!�f���>�̾��@�V��b��F���=lͿ`   `   *A��ޖ��c�h�p�>��Q���Ӿ廑��~>���s���#_�����Rx����#_�s������~>�廑���Ӿ�Q�p�>�c�h�ޖ��`   `   ��+��q%����������+�����G�Z�������H�9_��䆼��Q��䆼9_���H�����Z���G�+�������������q%�`   `   ��Ҿ�˾{����R�� 7w��-:��`�ֶ���q����Q�μ����^u������Q�μ�����q�ֶ��`��-:� 7w��R��{����˾`   `   ]�|���t��]^�{J>�� ��/���y����A�������h�X�޼�h��������A�y�������/�� �{J>��]^���t�`   `   ~�����p��Z���뽽�͚���}�w?X�E�w]A�ٟE���K��;N���K�ٟE�w]A�E�w?X���}��͚��뽽Z��p�����`   `   ����G󠽴���}��(�r��{_�YJ[��th�Ms��g5�������պ�~�����g5��Ms���th�YJ[��{_�(�r��}�����G�`   `   ,�2�G�0�T�,��+�e�3�b�K�Z�x���\ǽ�{�����_6�cm"�_6�����{���\ǽ�Z�x�b�K�e�3��+�T�,�G�0�`   `   �'����ża�ڼE����-�+�r�����&}���G��m�.����F��.����m���G��}��&����+�r���-�E��a�ڼ��ż`   `   zWe��n�������L��W�8��6���7��z��(������r־p�޾r־�����(���z��7��6��8��W��L������n��`   `   I\;�ul�C�ż�.�����k���F>�ߍ���������	��*+��(2��*+�	��������ߍ���F>��k������.�C�żul�`   `   ƘZ��*��[����p�Z�ӽ40�����zeξ:3���?��,l�I[���`��I[���,l���?�:3�zeξ����40�Z�ӽ��p�[���*��`   `   ����ż�2�$礽���ܤt��þ���{dT�n`�������ϿCڿ��Ͽ���n`��{dT�����þܤt����$礽�2��ż`   `   �fʼ���Rl���ٽ�A��j���>�W�L�F���B�п�aA��m'�aA��B�пF���W�L��>��j���A���ٽ�Rl���`   `   ����+���}|	���t�2Ѿ��+�I·��jͿ����C�'�l���|�'�l���C����jͿI·���+�2Ѿ��t�}|	����+�`   `   �"�w�P�C��̬%�䓾���e�T�@ث����pF�פ��O������O���פ��pF����@ث�e�T����䓾̬%�C��w�P�`   `   /�<�SDr�
�н�5>��<��t��>�y�kͿ!$�*C|��n��%��uW�%���n��*C|�!$�kͿ>�y�t���<���5>�
�нSDr�`   `   J�P��^��o���O��#��uV"��$�������:���������R&����������:�����$��uV"��#����O�o佪^��`   `   ��Z��t����r�W�1���J(�Ka���h���C�����s%���"�F�3��"�s%��������C��h�Ka���J(�1��r�W����t��`   `   \WY��n�����U�����K�$��s��H�-�;���������
��Q&��
��������-�;�H翄s��K�$�����U���뽠n��`   `   �HL�@����ݽM�G�5ٰ��
���~���Ͽ9%�S�|�陷��%��pO��%��陷�S�|�9%���Ͽ��~��
�5ٰ�M�G���ݽ@��`   `   �5���g��ƽ�$2�+s�������Z��Ӯ�S��T=G��ŉ�W����Q��W����ŉ�T=G�S���Ӯ���Z����+s���$2��ƽ��g�`   `   2���B�J֧�������A�ܾT-2��ڊ���Ͽ���^�C��l�8D|��l�^�C������Ͽ�ڊ�T-2�B�ܾ������J֧��B�`   `   ���H������|N��R�@K��p
���Q��n��Usѿv)��_�3V&��_�v)�Usѿ�n����Q�p
�@K���R�|N󽷹��H��`   `   ޫ�Q%�qtM��Ѻ�}!�f���>�̾��@�V��b��F���=lͿ z׿=lͿF����b��@�V���>�̾f���}!��Ѻ�qtM�Q%�`   `   �Rx����#_�s������~>�廑���Ӿ�Q�p�>�c�h�ޖ��*A��ޖ��c�h�p�>��Q���Ӿ廑��~>���s���#_����`   `   �.��5��㩼�a�e���$Mս�. �P�c��ؘ�>���q�澄� �	D��� �q��>����ؘ�P�c��. �$Mսe����a��㩼�5�`   `   <.��xL�U'���;�>�<��{��M�ӽ����C��Wu������㟾d���㟾�����Wu��C����N�ӽ�{��>�<��;�U'���xL�`   `   V����멼����>����>�H����չ�_�����-�R?�	�E�R?��-����_��չ���>�H����>㼳����멼`   `   H�!�y�C:��*��_�"�7�=���g��쎽����Fƽ�ؽ�L߽�ؽFƽ�����쎽��g�7�=�"��_��*�C:�z�`   `   �������W�����j���H��-�*�����3)��}<��OQ�]"a��g�]"a��OQ��}<��3)���*���-���H���j�W������`   `   V.�n������ý0�����p��*5�}�
��*㼊.̼ �Ƽ�yȼa ʼ�yȼ �Ƽ�.̼�*�}�
��*5���p�1����ý��n���`   `   �$[���S�qy>�\$ ����˹��倽�,)���Լg����*�ZJ���=߻ZJ����*�g����Լ�,)��倽˹����\$ �qy>���S�`   `   Qް�t���vᘾmi� G������Ľ^�v������	u����!����:��!�	u�������^�v���Ľ��� G�mi�vᘾt���`   `   '
�0��]���ž@Ҙ���\����4Ź��?Q�WǼ�����)�:�)�;�)�:����WǼ�?Q�4Ź������\�@Ҙ��ž]��0��`   `   U�U��(M�X�5�����K������Y��3��ɛ�y�G�j�O�ֺ�;;O�ֺF�j�y��ɛ��3��Y������K����X�5��(M�`   `   �	���癿������Y��#����[J��ZJ?�h�ݽM�f��=ɼ.����k�.����=ɼM�f�h�ݽZJ?�[J������#���Y������癿`   `   ��he��¿�L��mc�$��B�ξ>���m�R7���[�D�}����D�}��[�R7���m�>��B�ξ$��mc��L���¿he�`   `   Q{)�C" �2����ҿm旿GZN�cA�F����D?�A�нtQ�aLǼp��aLǼtQ�A�н�D?�F���cA�GZN�m旿��ҿ2��C" �`   `   \�h�}_Z�m�5�;t	��Z��[�����#�L�Ǿ�h�b �I���0��d��0�I���b ��h�L�Ǿ��#�[����Z��;t	�m�5�}_Z�`   `   4���}��1�d���(�]��旿��>�=��[1�����rG���(�3����(�rG�����[1��=�澾�>��旿]过�(�1�d��}��`   `   Z����o���-����@�U��%���E�Q�����b����#�a�����A�P\���A�a�����#�b������E�Q�%���U����@��-���o��`   `   v]��yӰ��}��{�I�������>�Y��"��Θ�Q+������P�|O��P�����Q+��Θ��"�>�Y�������{�I��}��yӰ�`   `   	����t��4D���%A���N���T;T�m� ������)�R���ܿR�3'!�ܿR�R����)�����m� �T;T�N������%A�4D���t��`   `   '(��5~��d-e�N})����ꙿ7�B�h�� ��ϯ�qyH�}��qyH��ϯ� ���h��7�B��ꙿ��N})�d-e�5~��`   `   `�h�-9Z���5��
��kÿ�9���)��Ѿ�xz��5�W����53����53�W����5��xz��Ѿ�)��9���kÿ�
���5�-9Z�`   `   ��(�7�������ӿ�뙿�S���F����S��C�z���� ���� �z����C󽇓S��F����S��뙿��ӿ���7��`   `   �C�x�߿¿
䚿_�f��x"�f�پ�o��b	*��Ľ�uU�0����0���uU��Ľb	*��o��f�پ�x"�_�f�
䚿¿x�߿`   `   Ͷ��K藿���e�Y�1�%����8񢾫�S��������� �﫩��r�﫩��� ���������S�8񢾐��1�%�e�Y����K藿`   `   5lP�`VH�_H2�
���f�E�� Xi�9e����Z���e�k�{#�e�k����Z���9e�Xi�E���f�
��_H2�`VH�`   `   	D��� �q��>����ؘ�P�c��. �$Mսe����a��㩼�5��.��5��㩼�a�e���$Mս�. �P�c��ؘ�>���q�澄� �`   `   d���㟾�����Wu��C����N�ӽ�{��>�<��;�U'���xL�<.��xL�U'���;�>�<��{��N�ӽ����C��Wu������㟾`   `   	�E�R?��-����`��չ���>�H����>㼳����멼V����멼����>����>�H����չ�`�����-�R?�`   `   �L߽�ؽFƽ�����쎽��g�7�=�"��_��*�C:�z�H�!�z�C:��*��_�"�7�=���g��쎽����Fƽ�ؽ`   `   �g�]"a��OQ��}<��3)���*���-���H���j�W�������������W�����j���H��-�*�����3)��}<��OQ�]"a�`   `   a ʼ�yȼ�Ƽ�.̼�*�}�
��*5���p�1����ý��n���V.�n������ý1�����p��*5�}�
��*㼊.̼ �Ƽ�yȼ`   `   �=߻[J����*�g����Լ�,)��倽˹����\$ �qy>���S��$[���S�qy>�\$ ����˹��倽�,)���Լg����*�[J��`   `   ���:��!�
u�������^�v���Ľ��� G�mi�vᘾt���Qް�t���vᘾmi� G������Ľ^�v������	u���!�`   `   �)�;�)�:����WǼ�?Q�4Ź������\�@Ҙ��ž]��0��'
�0��]���ž@Ҙ���\����4Ź��?Q�WǼ�����)�:`   `   �;;P�ֺG�j�y��ɛ��3��Y������K����X�5��(M�U�U��(M�X�5�����K������Y��3��ɛ�y�G�j�P�ֺ`   `   �k�.����=ɼM�f�h�ݽZJ?�[J������#���Y������癿�	���癿������Y��#����[J��ZJ?�h�ݽM�f��=ɼ.���`   `   ���D�}��[�R7���m�>��C�ξ$��mc��L���¿he���he��¿�L��mc�$��B�ξ>���m�R7���[�D�}�`   `   p��aLǼtQ�A�н�D?�F���cA�GZN�m旿��ҿ2��C" �Q{)�C" �2����ҿm旿GZN�cA�F����D?�A�нtQ�aLǼ`   `   �d��0�I���b ��h�L�Ǿ��#�[����Z��;t	�m�5�}_Z�\�h�}_Z�m�5�;t	��Z��[�����#�L�Ǿ�h�b �I���0�`   `   3����(�rG�����[1��=�澾�>��旿]过�(�1�d��}��4���}��1�d���(�]��旿��>�=��[1�����rG���(�`   `   P\���A�a�����#�b������E�Q�%���U����@��-���o��Z����o���-����@�U��%���E�Q�����b����#�a�����A�`   `   |O��P�����Q+��Θ��"�>�Y�������{�I��}��yӰ�v]��yӰ��}��{�I�������>�Y��"��Θ�Q+������P�`   `   3'!�ܿR�R����)�����m� �T;T�N������%A�4D���t��	����t��4D���%A���N���T;T�m� ������)�R���ܿR�`   `   |��qyH��ϯ� ���h��7�B��ꙿ��N})�d-e�5~��'(��5~��d-e�N})����ꙿ7�B�h�� ��ϯ�qyH�`   `   ���53�W����5��xz��Ѿ�)��9���kÿ�
���5�-9Z�`�h�-9Z���5��
��kÿ�9���)��Ѿ�xz��5�W����53�`   `   ��� �z����C󽇓S��F����S��뙿��ӿ���7����(�7�������ӿ�뙿�S���F����S��C�z���� �`   `   ��/���uU��Ľb	*��o��f�پ�x"�_�f�
䚿¿x�߿�C�x�߿¿
䚿_�f��x"�f�پ�o��b	*��Ľ�uU�/��`   `   �r���� ���������S�8񢾐��1�%�e�Y����K藿Ͷ��K藿���e�Y�1�%����8񢾫�S��������� ��`   `    {#�e�k����Z���9e�Xi�E���f�
��_H2�`VH�5lP�`VH�_H2�
���f�E��Xi�9e����Z���e�k�`   `   �\ ��⠻�FN�i�׼��B�i��M�p�)�֚b�{���sӨ����Q������sӨ�{���֚b�p�)�M�i����B�i�׼�FN��⠻`   `   Q��[DŻ��.��z��PW��Q�����&۽a.�<`5��-U�;+k�s�;+k��-U�<`5�a.��&۽����Q�PW��z����.�[DŻ`   `   F��SN���j�J���Ǽ&����D��I��U���f�ٽ�~���������~��f�ٽU����I����D�&���ǼJ����j��SN�`   `   ���Atܼ�vҼ��ȼsȼ� ټԲ��J����E��p���������᝽��������p���E�J��ղ��� ټsȼ��ȼ�vҼAtܼ`   `   �~\���U��pB�
�'����lc�ն̼��żs�Ѽу�ta��U�r��U�ta�у�t�Ѽ��żֶ̼lc����
�'��pB���U�`   `   I�Ľj���,�����)�b�i�'�!?�P���xl��<�3�)�C<&��~&�C<&�3�)��<�xl�P���!?�i�'�)�b����,��j���`   `   �$�������r8� >��]=���[1�9�Ѽ��O�e�����:��v;�;��v;���:f����O�9�Ѽ�[1�]=�� >��r8ｅ�����`   `   쐃�o�}��c��>��%�gpսt����k$�n�� ���/k�;Hn'<B~A<Hn'</k�; ���n���k$�t���gpս�%��>��c�o�}�`   `   /V˾��þX]�����݌b��r#�h�ٽ�Y���K�y�&���w;�3;<j�b<�3;<��w;y�&��K��Y��h�ٽ�r#�݌b����X]����þ`   `   N��<������=ؾ�����o��} ���Ľ�S��K��,�ۺ�<� I<�<,�ۺ�K���S���Ľ�} ��o������=ؾ���<��`   `   ��^���U�N=����CO��̨�k�a����1���sG�Ʃ%�0|y;�`<0|y;Ʃ%�sG�1������k�a��̨�CO����N=���U�`   `   ������T���V�S*!�����]��~<�ؽ��Y��_��9D��&;9D��_����Y�ؽ~<��]�����S*!��V��T�����`   `   yؿ%�Ϳ�M�����<�R�������p�p���������.�������.�������p�p�������<�R�����M��%�Ϳ`   `   �;��I@忙賿nY��g�4����W[���+������1������.�����1������+�W[�����g�4�nY���賿I@�;��`   `   M�-�$���<׿����}�R����˨�F�nnٽ{�Z���м�q����м{�Z�nnٽF��˨���}�R�����<׿��$�`   `   u�F� �:��9�J��:竿�h���D����zY����:Cz�j�����j��:Cz�����zY�D������h�:竿J���9� �:�`   `   XP���C��$�s���EP���Cp�e������'�b���������m��˼�m��������'�b�����e���Cp�EP��s����$���C�`   `   ��F��:��Z��~�ڠ��Ӿi��a�g6��3�_�c���H����Qռ���H��c��3�_�g6���a�Ӿi�ڠ���~��Z��:�`   `   z�-�u$��>�qؿ�D��n�U����a��BR��$�C�������gͼ���C����$�BR��a����n�U��D��qؿ�>�u$�`   `   o������忆ി�턿G�8�����x���{;�yGֽ��f� ���>׵� �����f�yGֽ�{;�x������G�8��턿�ി�忦��`   `   ,>׿�"Ϳ6Q���掿��U��3��_˾i�����&ٵ��CB�X�̼����X�̼�CB�&ٵ����i���_˾�3���U��掿6Q���"Ϳ`   `   ��������Wꃿ��V���#���뾂㠾;�P������ב�@��s��5QR�s��@���ב�����;�P��㠾��뾍�#���V�Wꃿ����`   `   !d[���R�L;�}��W�ﾰg��q�r�e���ý|\�Q]߼\�M���\�M�Q]߼|\��ýe��q�r��g��W��}��L;���R�`   `   �S����� ��s־L��+�y��.�k��
���1�SF������Ӄ����SF���1��
��k��.�+�y�L���s־� ����`   `   Q������sӨ�{���֚b�p�)�M�i����B�i�׼�FN��⠻�\ ��⠻�FN�i�׼��B�i��M�p�)�֚b�{���sӨ����`   `   s�;+k��-U�<`5�a.��&۽����Q�PW��z����.�\DŻQ��\DŻ��.��z��PW��Q�����&۽a.�<`5��-U�;+k�`   `   �����~��f�ٽU����I����D�&���ǼJ����j��SN�F��SN���j�J���Ǽ&����D��I��U���f�ٽ�~����`   `   �᝽��������p���E�J��ղ��� ټsȼ��ȼ�vҼAtܼ���Atܼ�vҼ��ȼsȼ� ټղ��J����E��p��������`   `   r��U�ta�҃�t�Ѽ��żֶ̼lc����
�'��pB���U��~\���U��pB�
�'����lc�ֶ̼��żt�Ѽу�ta��U�`   `   �~&�D<&�4�)��<�xl�Q���"?�i�'�*�b����,��k���I�Ľk���,�����)�b�i�'�!?�P���xl��<�4�)�D<&�`   `   �;��v;���:f����O�9�Ѽ�[1�]=�� >��r8ｅ������$�������r8� >��]=���[1�9�Ѽ��O�f�����:��v;`   `   B~A<Hn'<.k�; ���n���k$�t���gpս�%��>��c�o�}�쐃�o�}��c��>��%�gpսt����k$�n�� ���.k�;Hn'<`   `   j�b<�3;<��w;z�&��K��Y��h�ٽ�r#�݌b����X]����þ/V˾��þX]�����݌b��r#�h�ٽ�Y���K�z�&���w;�3;<`   `   � I<�<,�ۺ�K���S���Ľ�} ��o������=ؾ���<��N��<������=ؾ�����o��} ���Ľ�S��K��-�ۺ�<`   `   �`<0|y;Ʃ%�sG�1������k�a��̨�CO����N=���U���^���U�N=����CO��̨�k�a����1���sG�Ʃ%�0|y;`   `   �&;8D��_����Y�ؽ~<��]�����S*!��V��T�����������T���V�S*!�����]��~<�ؽ��Y��_��9D�`   `   ������.�������p�p�������<�R�����M��%�Ϳyؿ%�Ϳ�M�����<�R�������p�p���������.�`   `   ��.�����1������+�W[�����g�4�nY���賿I@�;���;��I@忙賿nY��g�4����W[���+������1����`   `   �q����м{�Z�nnٽF��˨���}�R�����<׿��$�M�-�$���<׿����}�R����˨�F�nnٽ{�Z���м`   `   ���j��:Cz�����zY�D������h�:竿J���9� �:�u�F� �:��9�J��:竿�h���D����zY����:Cz�j��`   `   �˼�m��������'�b�����e���Cp�EP��s����$���C�XP���C��$�s���EP���Cp�e������'�b���������m�`   `   Qռ���H��c��3�_�g6���a�Ӿi�ڠ���~��Z��:���F��:��Z��~�ڠ��Ӿi��a�g6��3�_�c���H����`   `   �gͼ���C����$�BR��a����n�U��D��qؿ�>�u$�z�-�u$��>�qؿ�D��n�U����a��BR��$�C������`   `   =׵� �����f�yGֽ�{;�x������G�8��턿�ി�忦��o������忆ി�턿G�8�����x���{;�yGֽ��f� ���`   `   ����W�̼�CB�&ٵ����i���_˾�3���U��掿6Q���"Ϳ,>׿�"Ϳ6Q���掿��U��3��_˾i�����&ٵ��CB�X�̼`   `   5QR�s��@���ב�����;�P��㠾��뾍�#���V�Wꃿ������������Wꃿ��V���#���뾂㠾;�P������ב�@��s��`   `   ��[�M�Q]߼|\��ýe��q�r��g��W��}��L;���R� d[���R�L;�}��W�ﾰg��q�r�e���ý|\�Q]߼[�M�`   `   �Ӄ����SF���1��
��k��.�+�y�L���s־� �����S����� ��s־L��+�y��.�k��
���1�SF�����`   `   �X;XA�:��T}p�Qm��8gU�W���[��Ǿ� �D���g�L��J.��L����g� �D�Ǿ�\��W���8gU�Rm��U}p���UA�:`   `   w��:we :V<�F�������i��uP�M��ǽMI��w��m!���&��m!�w�MI��ǽM���uP��i�����G��Y<�se :`   `   ������w���j����S���������7.�4�h�%ב�A���82��~zý82��A���&ב�4�h��7.����������S�j��x������`   `   �?~�طw���g�Q�W�QT���h��A��i�����-�C�/�>�B�6qI�>�B�C�/��-���i���A����h�QT�R�W���g�طw�`   `   ��ٜ
��M��ָϼ[s��OU~��L��:�S.E���b�����uݑ�nH��uݑ�������b�T.E��:��L�PU~�[s��׸ϼ�M��ٜ
�`   `   �E ���Jh�(�?������ɼ��y��R�0�^���7�ț:��v:���:��v:ě:��7�1�^��R���y���ɼ���)�?��Jh�E ��`   `   oR�'&ݽ/ƽ�����s{�.��nҼ>�D���:�;�y<��@<yPL<��@<�y<�:�;Ę�>�D��nҼ.��s{�����/ƽ'&ݽ`   `   H7�D�0�Z���D��̽z����4����5�ͻڅ�;�6Q<�]�<��<�]�<�6Q<م�;5�ͻ�����4�z���̽�D�Z��D�0�`   `   ���T���I�q�b�I�E��Kv��đ��)#�sY��WX:�A<'��<�<'��<�A<UX:sY���)#��đ�Kv�E��b�I�I�q�T���`   `   ��;�ƾ�T��𷓾�8e�vD%��۽A���L���`��;�<�< �<�<�<`��;�L��A����۽vD%��8e�𷓾�T���ƾ`   `   Z9��������s�Ͼ���wg�Z��"��W�G��}�:NxA<۵y<NxA<}�:�W�G�"��Z���wg���s�Ͼ�������`   `   ��H�}�@���*��{�Br׾����%�O��� ������ ����:��;��-<:��;��绶� ������ �%�O�����Br׾�{���*�}�@�`   `   ㊄���}�`�_�B6�	^
��Cž�&���Z%����c:������t9&g�;�t9�����c:����Z%��&���Cž	^
�B6�`�_���}�`   `   ����U}��{���.a�ht)�d�����G�H���|lr��l˼^zʻ]p��^zʻ�l˼|lr���G�H����d��ht)��.a�{��U}��`   `   �ƿY����ɤ���?�D�3_
��
��Mvg�h�ج������C������C���ج��h�Mvg��
��3_
�?�D����ɤ�Y���`   `   :�ݿ�=ӿ5䶿���*@X�"N�1�Ⱦ}�B��fУ�������������fУ�B��}�1�Ⱦ"N�*@X����5䶿�=ӿ`   `   
t�8ۿِ��¿��Ԍ_��[���ϾPI�����8�����-������cK�������-�8������PI����Ͼ�[�Ԍ_�¿��ِ��8ۿ`   `   
�ݿhIӿ�����hIY�Ւ���˾Q���R�ӹ���<1�M3���`�M3���<1�ӹ���R�Q����˾Ւ�hIY������hIӿ`   `   ��ƿב��d��l��� �F�c��+���q��/�~����(��ԣ��Y��ԣ���(�~���/��q�+��c�� �F�l���d��ב��`   `   ����zW��������b�/�+�����Ŧ��V���8$��YM����9��YM�8$�����V��Ŧ����/�+���b�����zW��`   `   ��r}�&�_�;N7�����˾e����w5�\-ݽ�x���")^����")^����x�\-ݽ�w5�e����˾���;N7�&�_�r}�`   `   ��F��=?��G*�),��o۾�Π���^�S���5��,�C��<������7������<��,�C��5��S����^��Π��o۾),��G*��=?�`   `   ���c
�`'����Ͼ�V��X�q�w�(��:ݽ���2��|L|�'2��_M�'2��|L|�2������:ݽw�(�X�q��V����Ͼ`'��c
�`   `   �Ǿ�6���S���U���h��;-����+�����<�M������F�Z';F����M�����<�+������;-��h��U���S���6��`   `   J.��L����g� �D�Ǿ�\��W���8gU�Rm��U}p���TA�:�X;TA�:��U}p�Rm��8gU�W���\��Ǿ� �D���g�L��`   `   ��&��m!�w�MI��ǽM���uP��i�����G��Y<�oe :t��:pe :Y<�F�������i��uP�M��ǽMI��w��m!�`   `   zý82��A���&ב�4�h��7.����������S�k��x������������x���j����S���������7.�4�h�&ב�A���82��`   `   6qI�?�B�C�/��-���i���A����h�QT�R�W���g�طw��?~�طw���g�R�W�QT���h��A��i�����-�C�/�?�B�`   `   oH��vݑ�������b�T.E��:��L�PU~�[s��׸ϼ�M��ٜ
���ٜ
��M��׸ϼ[s��PU~��L��:�T.E���b�����vݑ�`   `   ���:��v:��:��7�2�^��R���y���ɼ���)�?��Jh�E ���E ���Jh�)�?������ɼ��y��R�1�^���7���:��v:`   `   xPL<��@<�y<�:�;Ƙ�?�D��nҼ.��s{�����/ƽ(&ݽoR�(&ݽ/ƽ�����s{�.��nҼ>�D�Ř��:�;�y<��@<`   `   ��<�]�<�6Q<م�;5�ͻ�����4�{���̽�D�Z��D�0�H7�D�0�Z���D��̽z����4����5�ͻم�;�6Q<�]�<`   `   �<'��<�A<SX:sY���)#��đ�Lv�E��b�I�I�q�T������T���I�q�b�I�E��Lv��đ��)#�sY��SX:�A<'��<`   `    �<�<�<`��;�L��A����۽vD%��8e�𷓾�T���ƾ��;�ƾ�T��𷓾�8e�vD%��۽A���L���`��;�<�<`   `   ۵y<NxA<}�:�W�G�"��Z���wg���s�Ͼ�������Z9��������s�Ͼ���wg�Z��"��W�G��}�:NxA<`   `   ��-<;��;��绶� ������ �%�O�����Br׾�{���*�}�@���H�}�@���*��{�Br׾����%�O��� ������ ����:��;`   `   'g�;�t9�����c:����Z%��&���Cž	^
�B6�`�_���}�㊄���}�`�_�B6�	^
��Cž�&���Z%����c:������t9`   `   Rp��]zʻ�l˼|lr���F�H����d��ht)��.a�{��U}������U}��{���.a�ht)�d�����G�H���|lr��l˼^zʻ`   `   �����C���ج��h�Mvg��
��3_
�?�D����ɤ�Y����ƿY����ɤ���?�D�3_
��
��Mvg�h�ج������C�`   `   �������fУ�B��}�1�Ⱦ"N�*@X����5䶿�=ӿ:�ݿ�=ӿ5䶿���*@X�"N�1�Ⱦ}�B��fУ������`   `   �cK�������-�7������PI����Ͼ�[�Ԍ_�¿��ِ��8ۿ
t�8ۿِ��¿��Ԍ_��[���ϾPI�����8�����-�����`   `   �`�M3���<1�ӹ���R�Q����˾Ւ�hIY������hIӿ
�ݿhIӿ�����hIY�Ւ���˾Q���R�ӹ���<1�M3��`   `   �Y��ԣ���(�~���/��q�+��c�� �F�l���d��ב����ƿב��d��l��� �F�c��+���q��/�~����(��ԣ�`   `   ��9��YM�8$�����V��Ŧ����/�+���b�����zW������zW��������b�/�+�����Ŧ��V���8$��YM��`   `   ���!)^����x�[-ݽ�w5�e����˾���;N7�&�_�r}���r}�&�_�;N7�����˾e����w5�\-ݽ�x���")^�`   `   �7������<��,�C��5��S����^��Π��o۾),��G*��=?���F��=?��G*�),��o۾�Π���^�S���5��,�C��<�����`   `   WM�&2��|L|�1������:ݽw�(�X�q��V����Ͼ`'��c
����c
�`'����Ͼ�V��X�q�w�(��:ݽ���2��|L|�'2��`   `   [';F����M�����<�+������;-��h��U���S���6���Ǿ�6���S���U���h��;-����+�����<�M������F�`   `   �<���;,yT;h��Fzw�`D��.uJ�����ǽ(��I���#�y�(��#�I��(����ǽ��.uJ�aD��Gzw�h��)yT;���;`   `   N3�;�D�;4�;�&�B��k�����{�3��Lv��A������%̽(ӽ%̽�����A���Lv�{�3����k��D��7�&�3�;�D�;`   `   ��d;�gT;V�;uZ	:�{/����,#k��庼���3,��2N�fpe���m�fpe��2N�3,�����庼-#k�����{/�kZ	:T�;�gT;`   `   �:��8I����q��>�R�+�ͤX�lL���]��:U��Ƒ��#��$�ͼʥּ$�ͼ�#���Ƒ��:U��]�mL��ФX�U�+��>���q�8I��`   `   h��P~���6w��<�;���膻rX޺���i-?�2���F�����񓻫����F�5��r-?����wX޺�膻;���<��6w�P~��`   `   Mn#��z�s���ؼϬ��z�*�şd�:3�:��;�� <�,<��<�<��<�,<�� <��;73�:ǟd�z�*�Ϭ���ؼs���z�`   `   >�)����x�(KJ���M���e/�0�;����;jNH<��<���<J�<���<��<jNH<���;6�;�e/�M�����(KJ���x�)��`   `   �&����˽�2���A~��x+��g������j{;��K<�<�<L�<�U�<L�<�<�<��K<�j{;����g���x+��A~��2���˽��`   `   ��3��p-����j��|�ǽ�勽��+��"���PE�bB<iˎ<�[�<�r�<�[�<iˎ<bB<�PE��"����+��勽|�ǽj������p-�`   `   4���4�{��?b��=������ѽ�z���(���V�a�a;d�k<�8�<�{�<�8�<d�k<`�a;��V��(��z����ѽ����=��?b�4�{�`   `   (������Bw��}����L������ý@e�`Լ����T�<��<׾�<��<T�<����`Լ@e���ý�����L�}��Bw������`   `   �5��b/�eIҾ��/釾_�D��+����R�%��b�'7k;�Z<_��<�Z<'7k;�b�R�%�����+�_�D�/釾��eIҾb/�`   `   ��������h�޾/V���~y��v(��+ѽ�2e�1�¼��B�۲<�CI<۲<��B�1�¼�2e��+ѽ�v(��~y�/V��h�޾�����`   `   ˦@�N9�m1$�gN��Jо�_����K��������	����~w;u:<�~w;��	����������K��_���JоgN�m1$�N9�`   `   
^`��6W�C\>�,�F`�\X��$ri���i;��t�+�w${���)����;��)�w${�t�+�i;����$ri�\X��F`�,�C\>��6W�`   `   �v��Ql�V�P�\�*��o� ���kH~�$�!��(��r�E��4W����=:3W���r�E��(��$�!�kH~� ����o�\�*�V�P��Ql�`   `   A�~��s�s9W���/�z�����ǁ��O1(��ǽ�5T��6���ۻp{Ӻ�ۻ�6���5T��ǽO1(�ǁ�����z����/�s9W��s�`   `   �v�+al���P�2 +��'��Y���(��&�2sƽ��U�N��?) �y07�?) �N����U�2sƽ&��(���Y���'�2 +���P�+al�`   `   "A`�C;W�}�>��������p�Ĭ�l��� 3J��Ϸ�
'����3�
'���Ϸ� 3J�l���Ĭ��p������}�>�C;W�`   `   tF@���8�
~$��C��Ӿn�����U�;�
�@����P3��E������>ɺ����E���P3�@���;�
���U�n����Ӿ�C�
~$���8�`   `   {0�Og����	{�0���0y����3�)��0������v�H�S�h�:G�S���v����0��)���3�0y��0���	{����Og�`   `   ����	�+vѾ��)Њ��N�����亽X2]�)�༝/"�ٴO�Q;M�O��/"�)��X2]��亽����N�)Њ���+vѾ�	�`   `   Lj���_��Q���߇��?�P�:���iٽ�<���!�����0���U;m˾;�U;�0������!��<���iٽ:��?�P�߇��Q����_��`   `   <�{��fs��`\��
;����:O޽1T��TnC�-�ּ�,��Y��k�;�|<k�;�Y���,�-�ּTnC�0T��:O޽����
;��`\��fs�`   `   y�(��#�I��(����ǽ��.uJ�aD��Gzw�h��)yT;���;�<���;)yT;h��Gzw�aD��.uJ�����ǽ(��I���#�`   `   (ӽ%̽�����A���Lv�{�3����k��D��9�&�3�;�D�;M3�;�D�;3�;3�&�D��k�����{�3��Lv��A������%̽`   `   ��m�fpe��2N�3,�����庼-#k�����{/�jZ	:S�;�gT;��d;�gT;S�;kZ	:�{/����-#k��庼���3,��2N�fpe�`   `   ʥּ$�ͼ�#���Ƒ��:U��]�mL��ФX�U�+���>���q�9I���:��9I����q���>�U�+�ФX�mL���]��:U��Ƒ��#��$�ͼ`   `   񓻫����F�6��s-?����xX޺�膻;���<��6w�P~��h��P~���6w��<�;���膻wX޺���r-?�6���F�����`   `   �<��<�,<�� <��;63�:ǟd�z�*�Ϭ���ؼs���z�Mn#��z�s���ؼϬ��z�*�ǟd�73�:��;�� <�,<��<`   `   J�<���<��<jNH<���;7�;�e/�M�����)KJ���x�)��>�)����x�)KJ���M���e/�7�;����;jNH<��<���<`   `   �U�<L�<�<�<��K<�j{;����g���x+��A~��2���˽�㽛&����˽�2���A~��x+��g������j{;��K<�<�<L�<`   `   �r�<�[�<iˎ<bB<�PE��"����+��勽|�ǽj������p-���3��p-����j��|�ǽ�勽��+��"���PE�bB<iˎ<�[�<`   `   �{�<�8�<d�k<a�a;��V��(��z����ѽ����=��?b�4�{�4���4�{��?b��=������ѽ�z���(���V�`�a;c�k<�8�<`   `   ׾�<��<T�<����`Լ@e���ý�����L�}��Bw������(������Bw��}����L������ý@e�`Լ����T�<��<`   `   _��<�Z<(7k;�b�R�%�����+�`�D�/釾��eIҾb/��5��b/�eIҾ��/釾`�D��+����R�%��b�'7k;�Z<`   `   �CI<ܲ<��B�0�¼�2e��+ѽ�v(��~y�/V��h�޾�������������h�޾/V���~y��v(��+ѽ�2e�1�¼��B�۲<`   `   v:<�~w;��	����������K��_���JоgN�m1$�N9�˦@�N9�m1$�gN��Jо�_����K��������	����~w;`   `   ���;��)�w${�t�+�i;����$ri�\X��F`�,�C\>��6W�
^`��6W�C\>�,�F`�\X��$ri���i;��t�+�w${���)�`   `   ��=:2W���r�E��(��$�!�kH~� ����o�\�*�V�P��Ql��v��Ql�V�P�\�*��o� ���kH~�$�!��(��r�E��3W��`   `   k{Ӻ�ۻ�6���5T��ǽO1(�ǁ�����z����/�s9W��s�A�~��s�s9W���/�z�����ǁ��O1(��ǽ�5T��6���ۻ`   `   v07�?) �N����U�2sƽ&��(���Y���'�2 +���P�+al��v�+al���P�2 +��'��Y���(��&�2sƽ��U�N��?) �`   `   ��3�	'���Ϸ� 3J�l���Ĭ��p������}�>�C;W�"A`�C;W�}�>��������p�Ĭ�l��� 3J��Ϸ�
'��`   `   �>ɺ����E���P3�@���;�
���U�n����Ӿ�C�
~$���8�tF@���8�
~$��C��Ӿn�����U�;�
�@����P3��E�����`   `   q�:D�S���v����0��(���3�0y��0���	{����Og�{0�Og����	{�0���0y����3�)��0������v�F�S�`   `   Q;!�O��/"�)��X2]��亽����N�)Њ���+vѾ�	龙���	�+vѾ��)Њ��N�����亽X2]�)�༝/"��O�`   `   n˾;�U;�0����� �!��<���iٽ:��?�P�߇��Q����_��Lj���_��Q���߇��?�P�:���iٽ�<���!�����0���U;`   `   �|< k�;X���,�-�ּSnC�0T��:O޽����
;��`\��fs�<�{��fs��`\��
;����:O޽1T��TnC�-�ּ�,�_Y��k�;`   `   )�\<��M<c�<�;��&�L���˼�!��b������ޫ�vL��o�ĽwL���ޫ������b��!���˼L���&��;c�<��M<`   `   �P<|iG<�,<J^�;��>;nG^���:��2��g����t)�K�L�|�d�mtm�|�d�K�L��t)�g����2����:�rG^���>;I^�;�,<|iG<`   `   �U"<c�<�c<&�<X@�;'-6;�ʺ���1�U�<����Ǽ���wB�����Ǽ<���1�U�����ʺ$-6;W@�;&�<�c<c�<`   `   gF�;�B�;�;��;� �; �;y�;�-;G�� H�?n��0���Y	�0���@n��H�UG���-;y�;�;� �;��;�;�B�;`   `   �F������K�%�邶L�6;&��;
��;��<�$< f <�U�;���;���;���;�U�; f <�$<��<	��;%��;J�6;5삶L�%�����`   `   2���|d���p��1"�m~����:�;�#<�dP<X�l<� |<���<$��<���<� |<X�l<�dP<�#<�;��:m~�� 2"��p�|d��`   `   �� �}o���~�˼�҂����Ș�:�X<8�`<��<G
�<��<Q��<��<G
�<��<8�`<�X<Ƙ�:��⻠҂�~�˼��}o�`   `   gy������6i���;��������u�5a;!�?<���<;��<NU�<M�<NU�<;��<���<!�?<5a;u����������;��6i����`   `   '?սqiͽR��Ӗ�\�a����ne��r����$�;=_�<�=�<u��<[{�<u��<�=�<=_�<�$�;r���ne�����\�a�Ӗ�R��qiͽ`   `   ������!�\=߽p&��7zm�����Hv�1�9a�?<��<�Y�<���<�Y�<��<a�?<1�9�Hv����7zm�p&��\=߽�!����`   `   �4V���N���9��i��!�N����{Z�g�����%�;v��<Yc�<��<Yc�<v��<�%�;��g�传{Z�N����!�i���9���N�`   `   !s���}��Xu�4|M�y< ��f�-���z-������Vj�:�@<��<jǨ<��<:�@<hVj������z-�-���f�y< �4|M�Xu��}��`   `   ����:Q��f����p��`&J�J����ĽCk��u伛�ݻ�/�;עv<s#�<עv<�/�;��ݻ�u�Ck���ĽJ��`&J��p��f���:Q��`   `   �o׾�Ͼ����k��X�r�A�0��;�qߒ����_OZ�D2+;,�=<�-m<,�=<D2+;_OZ����qߒ��;�A�0�X�r��k������Ͼ`   `   �%�� վU����w��s*J��	�?���x<�0'��Yú�H	<|M=<�H	<Yú0'��x<�?����	�s*J��w��U���� վ�`   `   l�In�2h�[����6����[���c��1�T��ʿ������c�;[�<�c�;�����ʿ�1�T�c������[��6��[���2h�In�`   `   �K
�](�?Xƾ����7�b�r�˧Ž��a�`�Լ�L�:�z;��;:�z;�L�`�Լ��a�˧Žr�7�b������Xƾ?�](�`   `   Gk��x����Ic��20���^�T����ýha��sؼ�����~:;�U�;�~:;�����sؼha���ýT���^�20��Ic����群x�`   `   �����o}վh���";��<�N�����`����S��_˼���R:;��;�R:;�黜_˼��S��`�����<�N�";��h���o}վ��`   `   q�־�cϾ�x��򷜾?w���6�U���Uâ�C�:�����P���<w;���;�<w;�P�����C�:�Uâ�U�����6�?w�򷜾�x���cϾ`   `   X���b���1���;���<�N����\ս�+��*�����i$���;u�<��;�i$����*��+��\ս���<�N�;���1���b���`   `   ӫ��f	���9t���N��_$�����?���"U���漽�0�^�i:e5�;U�<f5�;_�i:��0�����"U��?������_$���N��9t�f	��`   `   �Q��8J�A17��}��=��Ps��{������|g��7T�;��<��<<��<8T�;|g�������{�Ps���=���}�A17��8J�`   `   �:��k�z��rNܽ�g��[��7�*�
�ļ3#�\��9���;��=<�yS<��=<���;_��93#�	�ļ7�*�[���g��rNܽz���k�`   `   p�ĽwL���ޫ������b��!���˼L���&��;c�<��M<)�\<��M<c�<�;��&�L���˼�!��b������ޫ�wL��`   `   mtm�|�d�K�L��t)�g����2����:�rG^���>;I^�;�,<{iG<�P<{iG<�,<I^�;��>;rG^���:��2��g����t)�K�L�|�d�`   `   wB�����Ǽ<���1�U�����ʺ$-6;W@�;&�<�c<c�<�U"<c�<�c<&�<W@�;$-6;�ʺ���1�U�<����Ǽ���`   `   Z	�1���@n��H�YG���-;y�;�;� �;��;�;�B�;fF�;�B�;�;��;� �;�;y�;�-;QG��H�@n��1���`   `   ���;���;�U�; f <�$<��<	��;%��;J�6;z킶M�%������F������M�%�*킶J�6;%��;	��;��<�$< f <�U�;���;`   `   $��<���<� |<X�l<�dP<�#<�;��:n~�� 2"��p�|d��2���|d���p� 2"�n~����:�;�#<�dP<X�l<� |<���<`   `   Q��<��<G
�<��<8�`<�X<Ř�:��⻠҂�~�˼��}o��� �}o���~�˼�҂����Ř�:�X<8�`<��<G
�<��<`   `   M�<NU�<;��<���<!�?<5a;u����������;��6i����gy������6i���;��������u�5a;!�?<���<;��<NU�<`   `   [{�<u��<�=�<=_�<�$�;r���ne�����\�a�Ӗ�R��qiͽ'?սqiͽR��Ӗ�\�a����ne��s����$�;=_�<�=�<u��<`   `   ���<�Y�<��<a�?<1�9�Hv����7zm�p&��\=߽�!����������!�\=߽p&��7zm�����Hv�1�9a�?<��<�Y�<`   `   ��<Yc�<w��<�%�;��g�传{Z�N����!�i���9���N��4V���N���9��i��!�N����{Z�g�����%�;v��<Yc�<`   `   kǨ<��<:�@<XUj������z-�-���f�y< �4|M�Xu��}��!s���}��Xu�4|M�y< ��f�-���z-������Vj�:�@<��<`   `   s#�<עv<�/�;��ݻ�u�Ck���ĽJ��`&J��p��f���:Q������:Q��f����p��`&J�J����ĽCk��u伛�ݻ�/�;עv<`   `   �-m<-�=<F2+;_OZ����qߒ��;�A�0�X�r��k������Ͼ�o׾�Ͼ����k��X�r�A�0��;�qߒ����_OZ�D2+;,�=<`   `   |M=<�H	<Yú0'��x<�?����	�s*J��w��U���� վ%�� վU����w��s*J��	�?���x<�0'��Yú�H	<`   `   \�<�c�;�����ʿ�1�T�c������[��6��[���2h�In�l�In�2h�[����6����[���c��1�T��ʿ������c�;`   `   ��;=�z;�L�`�Լ��a�˧Žr�7�b������Xƾ?�](��K
�](�?Xƾ����7�b�r�˧Ž��a�`�Լ�L�<�z;`   `   �U�;�~:;�����sؼha���ýT���^�20��Ic����群x�Gk��x����Ic��20���^�T����ýha��sؼ�����~:;`   `   ��;�R:;�黛_˼��S��`�����<�N�!;��h���o}վ�������o}վh���";��<�N�����`����S��_˼���R:;`   `   ���;�<w;�P�����C�:�Uâ�T�����6�?w�򷜾�x���cϾq�־�cϾ�x��򷜾?w���6�U���Uâ�C�:�����P���<w;`   `   v�<��;�i$����*��+��\ս���<�N�;���1���b���X���b���1���;���<�N����\ս�+��*�����i$���;`   `   U�<g5�;l�i:��0�����"U��?������_$���N��9t�f	��ӫ��f	���9t���N��_$�����?���"U���漽�0�a�i:f5�;`   `   ��<<��<9T�;zg�������{�Ps���=���}�A17��8J��Q��8J�A17��}��=��Ps��{������|g��8T�;��<`   `   �yS<��=<���;y��92#�	�ļ7�*�[���g��rNܽz���k��:��k�z��rNܽ�g��[��7�*�
�ļ3#�^��9���;��=<`   `   ?��<i�<��t<4A<d�;;�:{ֻ�z�JOʼ�o
�*��W?���F��W?�*��o
�KOʼ�z�{ֻ3�:d�;4A<��t<h�<`   `   ��<h�<��|<��]<m/<��;���:��w��Q#��(��4���ɼ�Ӽ�ɼ4���(���Q#���w����:��;m/<��]<��|<h�<`   `   )*v<?�t<;:o<��c<�P<ݰ1<D�<��;U��:���Ϯ��e������e���Ϯ���O��:��;C�<ݰ1<�P<��c<::o<?�t<`   `   ��;<�q><x�D<��L<��R< �R<v!J<W8<,'<��<m��;�֭;y�;�֭;l��;��<,'<W8<u!J< �R<��R<��L<w�D<�q><`   `   �w�;�;�;���;�<4�1<��O<�f<St<�Rx<X�u<�vp<܈k<��i<ۈk<�vp<X�u<�Rx<St<�f<��O<3�1<�<���;�;�;`   `   /�S�T.#�:�͹�J3;+�;=&<n�\<	G�<�$�<	w�<�y�<{o�<>O�<{o�<�y�<	w�<�$�<	G�<n�\<=&<+�;�J3;A�͹T.#�`   `   ���ߩn�#�9�aջ�4P�
ܦ;v�,<��x<���<t��<ܪ�<���<�
�<���<ܪ�<t��<���<��x<v�,<	ܦ;�4P�aջ#�9�ߩn�`   `   Z6�������ּ����ir5��O*�/�;c�F<� �<�:�<���<Y^�<�v�<Y^�<���<�:�<� �<c�F<.�;�O*�ir5�������ּ����`   `   �_^�v�T��:��D�v�ɼA0U�����d�;D�p<�i�<���< ��<�E�< ��<���<�i�<D�p<�d�;���A0U�v�ɼ�D��:�v�T�`   `   F����>��d���h��%*���ռ.K@���:��*<=��<�n�<���< t�<���<�n�<=��<��*<��:.K@���ռ�%*��h�d���>��`   `   Lb轔��Ƚ����{��)�H�����r�;�+j<\�<+��<�R�<+��<\�<�+j<�r�;��H���)��{�����Ƚ��`   `   �C�.�������ݽ� ��zo�e��铅��щ��'<G��<�B�<���<�B�<G��<�'<�щ�蓅�e��zo�� ����ݽ���.��`   `   �I@��9��'�����ٽݙ��l�F��м�����;Dq<DO�<�گ<DO�<Dq<��;����мl�F�ݙ����ٽ���'��9�`   `   ��e���]���G��'��	�ur���fx������\�B��:K?<Ԏ<I'�<Ԏ<K?<C��:��\�����fx�ur���	��'���G���]�`   `   ]����e|��4c�b�>���y�ٽz��w�)�N��OM��<Gy<�e�<Gy<�<NM�N��w�)�z��y�ٽ��b�>��4c��e|�`   `   T^���y����u���N�3"�E;����fH?�����N������;�aZ<��}<�aZ<���;N�������fH?����E;�3"���N���u��y��`   `   �#��f"��cl|��bT��'��:��6 ��V�I�0�ɼ̏޻��;&RC<�pg<&RC<��;̏޻/�ɼV�I�6 ���:���'��bT�cl|�f"��`   `   �]�������%v�hO���#����簣�� H�˼�ﻴ��;j�5<�KY<j�5<���;��˼� H�簣������#�hO��%v�����`   `   u����q|���c��Y@�<���)�8�����:�GG����Ի��;��2< LT<��2<��;��ԻGG����:�8����)�<���Y@���c��q|�`   `   �0e���]��DH�f)�����Ž��� �"�~N���"���ӵ;��9<'|X<��9<�ӵ;�"��~N�� �"������Ž��f)��DH���]�`   `   <�>�ި8��'�����1ཋ���^�֥���n���кg�;�QI<"qd<�QI<g�;��к��n�֥��^�����1�����'�ި8�`   `   �����X)���߽�˰�-����*��M���6�&R�:�<�n^<ADu<�n^<�<'R�:�6��M����*�-���˰���߽X)����`   `   �L��ٽ.Žc5��})����:� �v1o�ؒH��F�;�<<I�t<ꍃ<I�t<�<<�F�;ؒH�v1o� ��:�})��c5��.Ž�ٽ`   `   �������ez����c���.�����$���`̻-�!;:�<jH]<�܃<�<�܃<jH]<:�<-�!;�`̻�$������.���c�ez������`   `   ��F��W?�*��o
�KOʼ�z�{ֻ3�:d�;4A<��t<h�<?��<h�<��t<4A<d�;4�:{ֻ�z�KOʼ�o
�*��W?�`   `   �Ӽ�ɼ4���(���Q#���w����:��;m/<��]<��|<g�<��<g�<��|<��]<m/<��;���:��w��Q#��(��4���ɼ`   `   ����e���Ϯ���O��:��;C�<ݰ1<�P<��c<::o<>�t<)*v<>�t<::o<��c<�P<ݰ1<C�<��;O��:���Ϯ��e��`   `   x�;�֭;l��;��<,'<W8<u!J< �R<��R<��L<w�D<�q><��;<�q><w�D<��L<��R< �R<u!J<W8<,'<��<l��;�֭;`   `   ��i<ۈk<�vp<X�u<�Rx<St<�f<��O<3�1<�<���;�;�;�w�;�;�;���;�<3�1<��O<�f<St<�Rx<X�u<�vp<ۈk<`   `   >O�<{o�<�y�<	w�<�$�<	G�<n�\<<&<+�;�J3;H�͹U.#�0�S�U.#�I�͹�J3;+�;<&<n�\<	G�<�$�<	w�<�y�<{o�<`   `   �
�<���<ܪ�<t��<���<��x<v�,<	ܦ;�4P�aջ$�9�ߩn����ߩn�$�9�aջ�4P�	ܦ;u�,<��x<���<t��<ܪ�<���<`   `   �v�<Y^�<���<�:�<� �<c�F<.�;�O*�jr5�������ּ����Z6�������ּ����jr5��O*�.�;c�F<� �<�:�<���<Y^�<`   `   �E�< ��<���<�i�<D�p<�d�;���A0U�v�ɼ�D��:�w�T��_^�w�T��:��D�v�ɼA0U�����d�;D�p<�i�<���< ��<`   `    t�<���<�n�<=��<��*<��:.K@���ռ�%*��h�d���>��F����>��d���h��%*���ռ/K@���:��*<=��<�n�<���<`   `   �R�<+��<\�<�+j<�r�;��H���)��{�����Ƚ��Lb轔��Ƚ����{��)�H�����r�;�+j<\�<+��<`   `   ���<�B�<G��<�'<�щ�蓅�e��zo�� ����ݽ���.���C�.�������ݽ� ��zo�e��铅��щ��'<G��<�B�<`   `   �گ<DO�<Dq<��;����мl�F�ݙ����ٽ���'��9��I@��9��'�����ٽݙ��l�F��м�����;Dq<DO�<`   `   I'�<	Ԏ<�K?<F��:��\�����fx�ur���	��'���G���]���e���]���G��'��	�ur���fx������\�B��:K?<Ԏ<`   `   �e�<Gy<�<LM�M��w�)�z��y�ٽ��b�>��4c��e|�]����e|��4c�b�>���y�ٽz��w�)�N��NM��<Gy<`   `   ��}<�aZ<���;M�������fH?����E;�3"���N���u��y��T^���y����u���N�3"�E;����fH?�����N������;�aZ<`   `   �pg<'RC<��;ʏ޻/�ɼV�I�6 ���:���'��bT�cl|�f"���#��f"��cl|��bT��'��:��6 ��V�I�0�ɼ̏޻��;'RC<`   `   �KY<j�5<���;��˼� H�簣������#�hO��%v������]�������%v�hO���#����簣�� H�˼�ﻴ��;j�5<`   `   LT<��2<��;��ԻGG����:�8����)�<���Y@���c��q|�u����q|���c��Y@�<���)�8�����:�GG����Ի��;��2<`   `   '|X<��9<�ӵ;�"��~N�� �"������Ž��f)��DH���]��0e���]��DH�f)�����Ž��� �"�~N���"���ӵ;��9<`   `   "qd<�QI<g�;y�к��n�֥��^�����1�����'�ި8�<�>�ި8��'�����1ཋ���^�֥���n���кg�;�QI<`   `   BDu<�n^<�<-R�:�6��M����*�-���˰���߽X)���������X)���߽�˰�-����*��M���6�&R�:�<�n^<`   `   ꍃ<I�t< �<<�F�;ԒH�u1o���:�|)��b5��.Ž�ٽ�L��ٽ.Žc5��})����:� �v1o�ؒH��F�;�<<I�t<`   `   �<�܃<kH]<;�<0�!;�`̻�$������.���c�ez�������������ez����c���.�����$���`̻-�!;:�<jH]<�܃<`   `   ���<)Ƣ<5�<g�<�j<490<���; �:��x��0��V��ނ�.���ނ��V��0���x��:���;390<�j<g�<5�<)Ƣ<`   `   �(�<M��<ڨ�<l�<Kʆ<��i<X=<�P<%מ;���:Zⶺ�Z��{���Z�]ⶺ���:$מ;�P<X=<��i<Kʆ<k�<٨�<M��<`   `   2z�<��<Rј<��<[(�<Z�<�`|<��_<�?<<}<���;3�;���;}<<�?<��_<�`|<Z�<[(�<��<Qј<��<`   `   '�<'
�<ym�<<g��<�<�ْ< �<���<U�<��t<��j<3sg<�j<��t<U�<���< �<�ْ<�<g��<<ym�<'
�<`   `   �Y<h�]<�Qj<�3}<bm�<z˓<�#�<s��<a.�<���<�<ű�<�I�<ű�<�<���<a.�<s��<�#�<y˓<bm�<�3}<�Qj<h�]<`   `   ��<�c<�>!<�B<�h<��<E�<{�<�G�<݈�<���<�Y�<��<�Y�<���<݈�<�G�<{�<D�<��<�h<�B<�>!<�c<`   `   iK:��:��c;Ĉ�;�#<!`<(+�<�E�<]�<�^�<���<�!�<���<�!�<���<�^�<]�<�E�<(+�<!`<�#<Ĉ�;��c;��:`   `   ��e� ��c��Jp�ud�;o�<5Rf<kȕ<Vű<{��<!7�<�~�<�0�<�~�<!7�<{��<Vű<kȕ<5Rf<o�<td�;Lp��c��e� �`   `   �n��2�������'p*�8v���N;��<��{<ף<;��<;9�<s��<�A�<s��<;9�<;��<ף<��{<��<��N;8v�'p*�����2���`   `   >�������Ｚ���QZ��r���K�;�;<Y��<��<�c�<��<f��<��<�c�<��<Y��<�;<�K�;�r���QZ������（��`   `   RY�AxP���6�5��R�ǼW0V��C!��$�;\�h<���<b�<�Q�<::�<�Q�<b�<���<\�h<�$�;�C!�W0V�R�Ǽ5����6�AxP�`   `   ��������	|�k�L��p�a��������:/�,<��<�ֳ<���<���<���<�ֳ<��</�,<���:���a���p�k�L��	|�����`   `   ։��0���8x��4��Z�G� �M���,�x�bU�;'�o<� �<Ya�<���<Ya�<� �<'�o<bU�;,�x�M��� �Z�G�4��8x��0���`   `   ,�04ٽ��½.ס���v��)���¼�`�)M;�E<��<:��<���<:��<��<�E<*M;�`���¼�)���v�.ס���½04ٽ`   `   �0 �	u���b޽���������G�o��F9V�w � �<zv�<揤<Z��<珤<zv�< �<�  �F9V�o����G���������b޽	u��`   `   G�
����𽗥ɽ�G���]�^S	��p��3��q� <�jr<��<���<��<�jr<r� <2���p��^S	��]��G����ɽ����`   `   �:��_	�$����ϽY����f���􋑼�$v�ݤ�;�`<ܝ�<�~�<ܝ�<�`<ޤ�;�$v�􋑼���f�Y�����Ͻ$���_	�`   `   ��
���'_��ʽ�
��A�a�@��?��E���I4�;ЦV<j�<(Ė<j�<ЦV<I4�;D���?��?��A�a��
���ʽ'_���`   `   ( �����>߽���)@��/�P� �C(���M����;�JU<Ԭ�<�Γ<Ԭ�<�JU<���;�M�C(���/�P�)@������>߽���`   `   �b���ؽ��ý2���C��4��߼a�R�	���X��;�H\<3y�<��<3y�<�H\<X��;���a�R��߼�4��C�2����ý��ؽ`   `   �����k������@��;�P��`��Ƭ�m����:1�<Ij<!�<�@�<!�<Ij<1�<���:m��Ƭ��`�;�P�@�������k��`   `   1e���U���z���O�Z����ӼÙe��r��'�;��5<Ǿ}<�ϓ<��<�ϓ<Ǿ}<��5<�'�;�r�Ùe���ӼZ����O��z��U��`   `   ��O�xH���1�I%�LԼ�[��qܻr��:m_<��X<�e�<9-�<���<9-�<�e�<��X<m_<s��:qܻ�[��LԼI%���1�xH�`   `   �������4߼E���h�JwݻfI9 <�;�T;<:~z<A�<���<wԣ<���<A�<:~z<�T;< <�;mI9Iwݻ�h�E��4߼����`   `   .���ނ��V��0���x��:���;390<�j<g�<5�<(Ƣ<���<(Ƣ<5�<g�<�j<390<���;�:��x��0��V��ނ�`   `   �{���Z�_ⶺ���:$מ;�P<X=<��i<Kʆ<k�<٨�<M��<�(�<M��<٨�<k�<Kʆ<��i<X=<�P<$מ;���:_ⶺ�Z�`   `   3�;���;}<<�?<��_<�`|<Z�<[(�<��<Qј<��<2z�<��<Qј<��<[(�<Z�<�`|<��_<�?<<}<���;`   `   3sg<�j<��t<U�<���< �<�ْ<�<g��<<ym�<'
�<'�<'
�<ym�<<g��<�<�ْ< �<���<U�<��t<�j<`   `   �I�<ű�<�<���<a.�<s��<�#�<y˓<bm�<�3}<�Qj<g�]<�Y<g�]<�Qj<�3}<bm�<y˓<�#�<s��<a.�<���<�<ű�<`   `   ��<�Y�<���<݈�<�G�<{�<D�<��<�h<�B<�>!<�c<��<�c<�>!<�B<�h<��<D�<{�<�G�<݈�<���<�Y�<`   `   ���<�!�<���<�^�<]�<�E�<(+�<!`<�#<È�;��c;��:dK:��:��c;È�;�#<!`<(+�<�E�<]�<�^�<���<�!�<`   `   �0�<�~�<!7�<{��<Vű<kȕ<5Rf<o�<td�;Op��c��f� ���f� ��c��Pp�td�;o�<5Rf<kȕ<Vű<{��<!7�<�~�<`   `   �A�<s��<;9�<;��<ף<��{<��<��N;8v�'p*�����2����n��2�������'p*�8v���N;��<��{<ף<;��<;9�<s��<`   `   f��<��<�c�<��<Y��<�;<�K�;�r���QZ������（��>�������Ｚ���QZ��r���K�;�;<Y��<��<�c�<��<`   `   ::�<�Q�<b�<���<\�h<�$�;�C!�W0V�R�Ǽ5����6�AxP�SY�AxP���6�5��R�ǼX0V��C!��$�;\�h<���<b�<�Q�<`   `   ���<���<�ֳ<��</�,<���:���a���p�k�L��	|�������������	|�k�L��p�a��������:/�,<��<�ֳ<���<`   `   ���<Ya�<� �<'�o<bU�;+�x�M��� �Z�G�4��8x��0���։��0���8x��4��Z�G� �M���-�x�aU�;'�o<� �<Ya�<`   `   ���<:��<��<�E<+M;�`���¼�)���v�.ס���½04ٽ,�04ٽ��½.ס���v��)���¼�`�)M;�E<��<:��<`   `   [��<珤<zv�<�<����E9V�o����G���������b޽	u���0 �	u���b޽���������G�o��F9V�� � �<zv�<珤<`   `   ���<��<�jr<r� <0���p��^S	��]��G����ɽ����G�
����𽗥ɽ�G���]�^S	��p��3��r� <�jr<��<`   `   �~�<ݝ�<�`<ߤ�;�$v�󋑼���f�Y�����Ͻ$���_	��:��_	�$����ϽY����f���􋑼�$v�ޤ�;�`<ݝ�<`   `   (Ė<k�<ЦV<J4�;C���?��?��A�a��
���ʽ'_�����
���'_��ʽ�
��A�a�@��?��D���I4�;ЦV<k�<`   `   �Γ<Ԭ�<�JU<���;�M�B(���/�P�)@������>߽���( �����>߽���)@��/�P� �C(���M����;�JU<Ԭ�<`   `   ��<3y�<�H\<Z��;���`�R��߼�4��C�2����ý��ؽ�b���ؽ��ý2���C��4��߼a�R�	���X��;�H\<3y�<`   `   �@�<!�<Jj<2�<���:m��Ƭ��`�;�P�@�������k�������k������@��;�P��`��Ƭ�m����:1�<Ij<!�<`   `   ��<�ϓ<Ǿ}<��5<�'�;�r�e���ӼY����O��z��U��1e���U���z���O�Z����ӼÙe��r��'�;��5<Ǿ}<�ϓ<`   `   ���<9-�<�e�<��X<n_<y��:oܻ�[��LԼI%���1�wH���O�xH���1�I%�LԼ�[��qܻq��:m_<��X<�e�<9-�<`   `   wԣ<���<A�<;~z<�T;<!<�;�I9Hwݻ�h�E��4߼�����������4߼E���h�JwݻeI9 <�;�T;<:~z<A�<���<`   `   ��<�h�<}��<h��<�G�< F�<�w<��M<O!<���;"u�;��k;qJ;��k;!u�;���;N!<��M<�w< F�<�G�<h��<}��<�h�<`   `   ���<�̴<�R�<X�<t��<�<.��<�d�<u�o<��S<�;<�n+<ý%<�n+<�;<��S<u�o<�d�<-��<�<t��<X�<�R�<�̴<`   `   Rְ<`��<l�<���<��<�ݪ<���<�[�<�~�<�[�<\-�<�4�<g�<�4�<\-�<�[�<�~�<�[�<���<�ݪ<��<���<l�<`��<`   `   ]X�<��<Bݩ<���<T�<!n�<�1�<�[�<��<$�<o��<�Y�<d{�<�Y�<n��<$�<��<�[�<�1�<!n�<T�<���<Bݩ<��<`   `   ���<�(�<�_�<g��<��<S�<$�<�r�<��<�/�<�X�<K-�<��<K-�<�X�<�/�<��<�r�<$�<S�<��<g��<�_�<�(�<`   `   �j�<�Ђ<���<ٓ<U�<�5�<Ձ�<���<]�<a�<1�<<��<�{�<<��<1�<a�<]�<���<Ձ�<�5�<U�<ٓ<���<�Ђ<`   `   H�@<CtG<��Z<�'x<+r�<b��<�}�<�$�<���<��<<��<���<$�<���<<��<��<���<�$�<�}�<b��<+r�<�'x<��Z<CtG<`   `   ���;�Y�;k�<}:7<�<f<���<��<�~�</�<б�<s�<+��<J�<+��<s�<б�</�<�~�<��<���<�<f<|:7<k�<�Y�;`   `    �S9�Gt:E;a��;��!<��a<Ē�<�w�<b~�<�U�<�</��<,�</��<�<�U�<b~�<�w�<Ē�<��a<��!<a��;E;�Gt:`   `   �.��b�ֻF���\D�7�l�;��<�Nm<Yǘ<�̴<w?�<]"�<E��<��<E��<]"�<w?�<�̴<Yǘ<�Nm<��<�l�;UD�7F���b�ֻ`   `   �@���w�L�A����������;M�2< v�<�<bH�<�<?�<_��<?�<�<bH�<�< v�<M�2<���;������L�A��w�`   `   S)ӼJ�Ǽ����ITl��4��iv8|��;��W<��<�f�<^�<z��<ܳ�<z��<^�<�f�<��<��W<|��;�iv8�4�HTl�����J�Ǽ`   `   ���3
�J��,��i�_�VQ����L;�'<�<r��<7��<	�<`��<	�<7��<r��<�<�'<��L;VQ��h�_�,��J���3
�`   `   ܣ5���-�������� ���|�P���;�9e<��<� �<� �<�^�<� �<� �<��<�9e<��;P��|�� ���������-�`   `   &�S��K�ؤ2���^�Ǽ$�_�n�m���;@|G<���<�<3[�<|	�<3[�<�<���<@|G<��;n�m�$�_�^�Ǽ��ؤ2��K�`   `   %sg�}S^��D�_����T��q��WcY;�D0<68�<��<>�<w5�<>�<��<68�<�D0<XcY;q��T�����_��D�}S^�`   `   �hn��,e��K�9s$����Y��Us�1�;Ѣ!<�	<��<�A�<�P�<�A�<��<�	<Ѣ!<2�;Us㻤Y�����9s$��K��,e�`   `   wvg���^�IE�������3Ό��߻c;9�<�)x<���<�˭<���<�˭<���<�)x<9�<c;�߻3Ό���缣��IE���^�`   `   vcS�N#K�i�3��-���м}+x�D��=�C;B$"<�4x<ؙ<�<V��<�<ؙ<�4x<B$"<>�C;D��}+x���м�-�i�3�N#K�`   `   ��4��U-���I��th���#@��H���;��0<��~<(��<�G�<�i�<�G�<(��<��~<��0<��;�H��#@�sh��I�����U-�`   `   �����E�S��,Vx�4�19ɻ�;9G<u��<�l�<�=�<���<�=�<�l�<u��<9G<ʻ�;�194��+Vx�S��E�`   `   O�ʼ����yP����s�J��ڋ�ʼ;L*<�'c<��<
�<<�t�<<
�<��<�'c<L*<ʼ;ً�J����s�yP������`   `   �o�~|`��a4�G_��B�|B;�Z <�G<:�<��<���<�˰<�ֳ<�˰<���<��<:�<�G<�Z <|B;�B�F_仇a4�~|`�`   `   ʇ���T���f$��	:���;<N
?<�t<��<��<yǬ<3��<K �<3��<yǬ<��<��<�t<N
?<<���;��	:�f$��T��`   `   qJ;��k;!u�;���;N!<��M<�w< F�<�G�<h��<|��<�h�<��<�h�<|��<h��<�G�< F�<�w<��M<N!<���;!u�;��k;`   `   ½%<�n+<�;<��S<u�o<�d�<-��<�<t��<X�<�R�<�̴<���<�̴<�R�<X�<t��<�<-��<�d�<u�o<��S<�;<�n+<`   `   g�<�4�<[-�<�[�<�~�<�[�<���<�ݪ<��<���<l�<`��<Rְ<`��<l�<���<��<�ݪ<���<�[�<�~�<�[�<[-�<�4�<`   `   d{�<�Y�<n��<$�<��<�[�<�1�<!n�<T�<���<Bݩ<��<]X�<��<Bݩ<���<T�<!n�<�1�<�[�<��<$�<n��<�Y�<`   `   ��<K-�<�X�<�/�<��<�r�<$�<S�<��<f��<�_�<�(�<���<�(�<�_�<f��<��<S�<#�<�r�<��<�/�<�X�<K-�<`   `   �{�<<��<1�<a�<]�<���<Ձ�<�5�<U�<ٓ<���<�Ђ<�j�<�Ђ<���<ٓ<U�<�5�<Ձ�<���<]�<a�<1�<<��<`   `   $�<���<<��<��<���<�$�<�}�<b��<+r�<�'x<��Z<BtG<H�@<BtG<��Z<�'x<+r�<b��<�}�<�$�<���<��<<��<���<`   `   J�<+��<s�<б�</�<�~�<��<���<�<f<|:7<j�<�Y�;���;�Y�;j�<|:7<�<f<���<��<�~�</�<ϱ�<s�<+��<`   `   ,�</��<�<�U�<b~�<�w�<Ē�<��a<��!<`��;E;�Gt:�S9�Gt:E;`��;��!<��a<Ē�<�w�<b~�<�U�<�</��<`   `   ��<E��<]"�<w?�<�̴<Yǘ<�Nm<��<�l�;D�7G���b�ֻ�.��b�ֻG����C�7�l�;��<�Nm<Yǘ<�̴<w?�<]"�<E��<`   `   _��<?�<�<bH�<�<!v�<M�2<���;������L�A���w��@����w�L�A����������;M�2< v�<�<bH�<�<?�<`   `   ܳ�<z��<^�<�f�<��<��W<|��;
jv8�4�ITl�����J�ǼS)ӼJ�Ǽ����ITl��4�iv8{��;��W<��<�f�<^�<z��<`   `   `��<	�<7��<r��<�<�'<��L;VQ��h�_�,��J���3
����3
�J��,��i�_�WQ����L;�'<�<r��<7��<	�<`   `   �^�<� �<� �<��<�9e<��;P��|�� ���������-�ܣ5���-�������� ���|�"P���;�9e<��<� �<� �<`   `   |	�<3[�<�<���<A|G<��;l�m�$�_�^�Ǽ��ؤ2��K�&�S��K�ؤ2���^�Ǽ$�_�o�m���;@|G<���<�<3[�<`   `   w5�<>�<��<68�<�D0<ZcY;q��T�����_��D�}S^�%sg�}S^��D�_����T��q��WcY;�D0<68�<��<>�<`   `   �P�<�A�<��<�	<Ѣ!<4�;Ts㻤Y�����8s$��K��,e��hn��,e��K�9s$����Y��Us�1�;Ѣ!<�	<��<�A�<`   `   ���<�˭<���<�)x<:�< c;�߻3Ό���缣��IE���^�wvg���^�IE�������3Ό��߻c;9�<�)x<���<�˭<`   `   V��<�<ؙ<�4x<C$"<A�C;C��|+x���м�-�h�3�N#K�ucS�N#K�i�3��-���м}+x�D��=�C;B$"<�4x<ؙ<�<`   `   �i�<�G�<(��<��~<��0<��;�H��#@�sh��H�����U-���4��U-���I��th���#@��H���;��0<��~<(��<�G�<`   `   ���<�=�<�l�<v��<�9G<˻�;�193��+Vx�S��E������E�S��,Vx�4�19ɻ�;9G<u��<�l�<�=�<`   `   �t�<<
�<��<�'c<M*<ͼ;֋�I����s�xP������O�ʼ����yP����s�J��ڋ�ʼ;L*<�'c<��<
�<<`   `   �ֳ<�˰<�<��<;�<�G<�Z <|B;�B�E_仆a4�~|`��o�~|`��a4�F_��B�|B;�Z <�G<:�<��<���<�˰<`   `   K �<3��<zǬ<��<��<�t<O
?<<���;��	:�f$��T��ʇ���T���f$��	:���;<N
?<�t<��<��<yǬ<3��<`   `   75�<�|�<ZT�<���<�÷<�4�<X�<��<���<��<v�<w�}<��y<w�}<v�<��<���<��<W�<�4�<�÷<���<ZT�<�|�<`   `   Ώ�<�A�<kU�<Pɿ<�t�<�$�<ﭵ<�*�<�<��<\��<�%�<1�<�%�<\��<��<�<�*�<ﭵ<�$�<�t�<Pɿ<kU�<�A�<`   `   C;�<jW�<٥�<u�<p4�<���<閿<�u�<1��<Xi�<'z�<�c�<6��<�c�<'z�<Xi�<1��<�u�<閿<���<p4�<u�<٥�<jW�<`   `   1��<J#�<H��<���<�~�<b��<�q�<?A�<�3�<U�<���<��<\K�<��<���<U�<�3�<?A�<�q�<b��<�~�<���<H��<J#�<`   `   ��<k�<�׷<��</��<���<��<���<)��<^�<�
�<5?�<J�<5?�<�
�<^�<)��<���<��<���</��<��<�׷<k�<`   `   /˨<�H�<Xq�<)��<��<�j�<3l�<�d�<��<�o�<���<���<�*�<���<���<�o�<��<�d�<3l�<�j�<��<)��<Xq�<�H�<`   `   �`�<xQ�<K�<�<�<"/�<G��<�k�<���<���<�-�<���<9��<���<9��<���<�-�<���<���<�k�<G��<"/�<�<�<K�<xQ�<`   `   �6�<��<j֎<���<́�<�<m�<��<���<w�<X�<w�<i�<w�<X�<w�<���<��<m�<�<́�<���<j֎<��<`   `   �;X<vy^<UQp<<]�<O�<���<6(�<v(�<Rb�<���<���<?(�<���<���<Rb�<v(�<6(�<���<O�<]�<<UQp<vy^<`   `   <r<>'$<�(:<]a[<뻁<q�<�M�<�T�<2;�<q��<Y��<���<J�<���<Y��<q��<2;�<�T�<�M�<q�<뻁<]a[<�(:<>'$<`   `   �*�;���;Xy�;%<̈U<+^�<~ߜ<���<���<�t�<�8�<B��<H��<B��<�8�<�t�<���<���<~ߜ<+^�<̈U<%<Xy�;���;`   `   �|:)��:�Lk;�d�;�+$<�`<Q.�<h��<�ֻ<o�<��<p?�<�u�<p?�<��<o�<�ֻ<h��<Q.�<�`<�+$<�d�;�Lk;)��:`   `   Te��K1����Xn@;M��;f8<<ez<.u�<���<;@�<o?�<1��<�W�<1��<o?�<;@�<���<.u�<=ez<f8<M��;Xn@;��깅K1�`   `   E���ۻv������Ɉ;�9<�4\< ��<��<�D�<b��<r�<@��<r�<b��<�D�<��<��<�4\<�9<Ɉ;���v����ۻ`   `   �n3��{#��l�n(J�cV�:_��;~VB<�Y�<P\�<��<q%�<{&�<��<{&�<q%�<��<P\�<�Y�<VB<_��;dV�:n(J��l��{#�`   `   �vW�x�F�s[������t9���;3:/<<�x<ޛ�<��<}
�<�m�<�{�<�m�<}
�<��<ޛ�<<�x<3:/<���;��t9���s[�x�F�`   `   i#d�ZVS��#�8鸻m��K��;��$<ߺn<��<_\�<���<�)�<�@�<�)�<���<_\�<��<ߺn<��$<K��;i��8鸻�#�ZVS�`   `   �W�KSG�Y�KE��!�,����;�$<��k<э�<�k�<*Y�<��<O��<��<*Y�<�k�<ҍ�<��k<�$<���;�,�JE��Y�KSG�`   `   ��2���#�Ʋ�2'g����:f�;�+-<!p<�Ǔ<�=�<�;�<O��<F��<O��<�;�<�=�<�Ǔ<!p<�+-<f�;���:2'g�Ʋ���#�`   `   ����xٻEB����l���R;M��;1?<3�z<�p�<iө<k�<�`�<_��<�`�<k�<iө<�p�<4�z<1?<M��;��R;��l�EB���xٻ`   `   8�K�&������;��;��<p�W<寅<�8�<��<r޷<Qؾ<�%�<Qؾ<r޷<��<�8�<寅<p�W<��< ��;��;���&�`   `   �1�:=�;�y;��;�<<E�E<�Lu<5�<8��<��<�h�<�A�<2�<�A�<�h�<��<8��<5�<�Lu<F�E<�<<��;�y;=�;`   `   ��;���;�<�n$<~I<7�o<\��<r(�<��<���<��<&_�<A��<&_�<��<���<��<r(�<\��<7�o<~I<�n$<�<���;`   `   <96<�y;<�sJ<�a<�S|< ��<�b�<홦<���<}��<�@�<a��<���<a��<�@�<~��<���<홦<�b�< ��<�S|<�a<�sJ<�y;<`   `   ��y<v�}<v�<��<���<��<W�<�4�<�÷<���<ZT�<�|�<65�<�|�<ZT�<���<�÷<�4�<W�<��<���<��<v�<v�}<`   `   1�<%�<\��<��<�<�*�<ﭵ<�$�<�t�<Pɿ<kU�<�A�<Ώ�<�A�<kU�<Pɿ<�t�<�$�<ﭵ<�*�<�<��<\��<%�<`   `   6��<�c�<'z�<Xi�<1��<�u�<閿<���<p4�<u�<٥�<jW�<C;�<jW�<٥�<u�<p4�<���<閿<�u�<1��<Xi�<'z�<�c�<`   `   \K�<��<���<U�<�3�<?A�<�q�<b��<�~�<���<H��<I#�<1��<I#�<H��<���<�~�<b��<�q�<?A�<�3�<U�<���<��<`   `   J�<5?�<�
�<^�<)��<���<��<���</��<��<�׷<k�<��<k�<�׷<��</��<���<��<���<)��<^�<�
�<5?�<`   `   �*�<���<���<�o�<��<�d�<3l�<�j�<��<)��<Xq�<�H�</˨<�H�<Xq�<)��<��<�j�<3l�<�d�<��<�o�<���<���<`   `   ���<8��<���<�-�<���<���<�k�<G��<"/�<�<�<K�<xQ�<�`�<xQ�<K�<�<�<"/�<G��<�k�<���<���<�-�<���<8��<`   `   i�<w�<X�<w�<���<��<m�<�<́�<���<j֎<��<�6�<��<j֎<���<́�<�<m�<��<���<w�<X�<w�<`   `   ?(�<���<���<Rb�<v(�<6(�<���<O�<]�<<UQp<vy^<�;X<vy^<UQp<<]�<O�<���<6(�<v(�<Rb�<���<���<`   `   J�<���<Y��<q��<2;�<�T�<�M�<q�<뻁<]a[<�(:<>'$<<r<>'$<�(:<]a[<뻁<q�<�M�<�T�<2;�<q��<Y��<���<`   `   H��<B��<�8�<�t�<���<���<~ߜ<+^�<̈U<%<Wy�;���;�*�;���;Wy�;%<̈U<+^�<~ߜ<���<���<�t�<�8�<B��<`   `   �u�<q?�<��<o�<�ֻ<h��<Q.�<�`<�+$<�d�;�Lk;(��:�|:'��:�Lk;�d�;�+$<�`<Q.�<h��<�ֻ<o�<��<p?�<`   `   �W�<1��<o?�<;@�<���<.u�<=ez<f8<M��;Xn@;��깆K1�Te��K1����Wn@;L��;f8<<ez<.u�<���<;@�<o?�<1��<`   `   @��<r�<b��<�D�<��<��<�4\<�9<Ɉ;���v����ۻE���ۻw������Ɉ;�9<�4\< ��<��<�D�<b��<r�<`   `   ��<{&�<r%�<��<P\�<�Y�<VB<`��;fV�:m(J��l��{#��n3��{#��l�o(J�bV�:_��;~VB<�Y�<P\�<��<q%�<{&�<`   `   �{�<�m�<}
�<��<ߛ�<=�x<3:/<���;�t9���s[�x�F��vW�x�F�s[������t9���;2:/<<�x<ޛ�<��<}
�<�m�<`   `   �@�<�)�<���<_\�<��<�n<��$<L��;\��8鸻�#�ZVS�i#d�ZVS��#�9鸻p��J��;��$<ߺn<��<_\�<���<�)�<`   `   O��<��<*Y�<�k�<ҍ�<��k<�$<���;��,�JE��Y�KSG��W�KSG�Y�KE��$�,����;�$<��k<э�<�k�<*Y�<��<`   `   F��<O��<�;�<�=�<�Ǔ<!p<�+-<h�;���:0'g�Ų���#���2���#�Ʋ�2'g����:f�;�+-<!p<�Ǔ<�=�<�;�<O��<`   `   _��<�`�<k�<jө<�p�<4�z<1?<O��;��R;��l�DB���xٻ����xٻEB����l���R;M��;1?<3�z<�p�<iө<k�<�`�<`   `   �%�<Qؾ<r޷<��<�8�<寅<q�W<��<!��;��;���&�7�K�&������; ��;��<p�W<寅<�8�<��<r޷<Qؾ<`   `   2�<�A�<�h�<��<8��<6�<�Lu<F�E<�<<��;�y;?�;�1�:>�;�y;��;�<<E�E<�Lu<5�<8��<��<�h�<�A�<`   `   A��<&_�<��<���<��<s(�<\��<8�o<~I<�n$<�<���;��;���;�<�n$<~I<7�o<\��<r(�<��<���<��<&_�<`   `   ���<a��<�@�<~��<���<홦<�b�< ��<�S|<�a<�sJ<�y;<=96<�y;<�sJ<�a<�S|< ��<�b�<홦<���<~��<�@�<a��<`   `   b��<(��<���<���<}��<Ť�<&4�<�F�<��<���<�P�<v��<I�<u��<�P�<���<��<�F�<&4�<Ť�<|��<���<���<(��<`   `   ��<o��<���<���<o{�<��<:�<���<\h�<q��<*A�<;�<<��<;�<*A�<q��<\h�<���<:�<��<o{�<���<���<o��<`   `   ���<E��<��<���<���<s��<�4�<�l�<�<�<	��<q2�<���<w��<���<p2�<	��<�<�<�l�<�4�<r��<���<���<��<E��<`   `   ��<�l�<@��<	��<���<���<y��<�f�<�g�<l��<�$�<�(�<�*�<�(�<�$�<l��<�g�<�f�<y��<���<���<	��<@��<�l�<`   `   ��<���<���<_�<���<��<�'�<��<s��<}P�<�,�<̘�<U��<̘�<�,�<}P�<s��<��<�'�<��<���<_�<���<���<`   `   ��<k��<*�<���<��<a��<��<���<,��<���<�s�<�>�<��<�>�<�s�<���<,��<���<��<`��<��<���<*�<k��<`   `   Qӻ<D޼<տ<�U�<���<���<8
�<���<+��<��<;"�<�S�<��<�S�<;"�<��<+��<���<8
�<���<���<�U�<տ<D޼<`   `   ��<d-�<0Ǹ<�7�<���<z��<��<޻�<.��<ӥ�<�]�<���<=��<���<�]�<ӥ�<.��<޻�<��<z��<���<�7�<0Ǹ<d-�<`   `   �<�o�<���<�O�<�@�<
��<���<@2�<�D�<��<�`�<�l�<��<�l�<�`�<��<�D�<@2�<���<
��<�@�<�O�<���<�o�<`   `   
�<_��<�ۤ<���< #�<�0�<��<]��<���<�S�<]�<���<���<���<]�<�S�<���<]��<��<�0�< #�<���<�ۤ<_��<`   `   � �<�C�<�_�<Ɨ�<���<��<���<���<kK�<���<o��<Ql�<�c�<Ql�<o��<���<kK�<���<���<��<���<Ɨ�<�_�<�C�<`   `   aH�<cŃ<���<Ԕ�<A{�<1�<�#�<F��<�R�<T��<�+�<�l�<؄�<�l�<�+�<T��<�R�<F��<�#�<1�<A{�<Ԕ�<���<cŃ<`   `   L�d<�Yj<��z<�h�<��<�i�<X �<�'�<��<�U�<�U�<���<'�<���<�U�<�U�<��<�'�<X �<�i�<��<�h�<��z<�Yj<`   `   TI<�dO<�Ha<�&|<~2�<#�<�O�<#��<�u�<��<p2�<��<Ni�<��<p2�<��<�u�<#��<�O�<#�<~2�<�&|<�Ha<�dO<`   `   ��2<�\9<�L<�Oi<�<z��<2A�<O��<?�<���< ��<<
�<�i�<=
�< ��<���<?�<O��<2A�<z��<�<�Oi<�L<�\9<`   `   ��#<k�*<��><�Y\<��<�<f�<�>�<^J�<�r�<���<���<�Q�<���<���<�r�<^J�<�>�<f�<�<��<�Y\<��><k�*<`   `   u�<�{%<;9<��V<�Oz<Ï<ԁ�<5�<�;�<Pd�<���<���<�F�<���<���<Pd�<�;�<5�<ԁ�<Ï<�Oz<��V<;9<�{%<`   `   R�#<�_*<t>=<��Y<h}{<D��<Ƒ�<���<J+�<���<���<�<8s�<�<���<���<J+�<���<Ƒ�<D��<i}{<��Y<t>=<�_*<`   `   �3<B9<�aJ<�Vd<���<~�<���<c��<�;�<�S�<���<D��<^ �<D��<���<�S�<�;�<c��<���<~�<���<�Vd<�aJ<B9<`   `   ��J<�2P<�X_<�v<终<�"�<��<�5�<x{�<��<�^�<���<��<���<�^�<��<x{�<�5�<��<�"�<终<�v<�X_<�2P<`   `   ��h<�hm<z<g��<V�<|'�<�ĩ<��<eɼ<u��<���<l��<���<l��<���<u��<eɼ<��<�ĩ<|'�<V�<g��<z<�hm<`   `   �D�<J	�<|�<]��<�ڜ<���<Hͯ<��<��<W��<���<��<���<��<���<W��<��<��<Hͯ<���<�ڜ<]��<|�<J	�<`   `   w�<�͗<枛<�]�<�F�<���<ً�<ν�<���<L�<\�<���<n��<���<\�<L�<���<ν�<ً�<���<�F�<�]�<枛<�͗<`   `   ���<&�<坪<;��<莳<���<�}�<���<K5�<���<��<mE�<d��<mE�<��<���<K5�<���<�}�<���<莳<;��<坪<&�<`   `   I�<u��<�P�<���<��<�F�<&4�<Ť�<|��<���<���<(��<b��<(��<���<���<|��<Ť�<&4�<�F�<��<���<�P�<u��<`   `   <��<;�<*A�<q��<\h�<���<:�<��<o{�<���<���<o��<��<o��<���<���<o{�<��<:�<���<\h�<q��<*A�<;�<`   `   w��<���<p2�<	��<�<�<�l�<�4�<r��<���<���<��<D��<���<D��<��<���<���<r��<�4�<�l�<�<�<	��<p2�<���<`   `   �*�<�(�<�$�<l��<�g�<�f�<y��<���<���<	��<@��<�l�<��<�l�<@��<	��<���<���<y��<�f�<�g�<l��<�$�<�(�<`   `   U��<̘�<�,�<}P�<s��<��<�'�<��<���<_�<���<���<��<���<���<_�<���<��<�'�<��<s��<}P�<�,�<̘�<`   `   ��<�>�<�s�<���<,��<���<��<`��<��<���<*�<k��<��<k��<*�<���<��<`��<��<���<,��<���<�s�<�>�<`   `   ��<�S�<;"�<��<+��<���<8
�<���<���<�U�<տ<D޼<Qӻ<D޼<տ<�U�<���<���<8
�<���<+��<��<;"�<�S�<`   `   =��<���<�]�<ӥ�<.��<޻�<��<z��<���<�7�<0Ǹ<d-�<��<d-�<0Ǹ<�7�<���<z��<��<޻�<.��<ӥ�<�]�<���<`   `   ��<�l�<�`�<��<�D�<@2�<���<
��<�@�<�O�<���<�o�<�<�o�<���<�O�<�@�<
��<���<@2�<�D�<��<�`�<�l�<`   `   ���<���<]�<�S�<���<]��<��<�0�< #�<���<�ۤ<_��<
�<_��<�ۤ<���<�"�<�0�<��<]��<���<�S�<]�<���<`   `   �c�<Ql�<o��<���<kK�<���<���<��<���<Ɨ�<�_�<�C�<� �<�C�<�_�<ŗ�<���<��<���<���<kK�<���<o��<Ql�<`   `   ؄�<�l�<�+�<T��<�R�<G��<�#�<1�<A{�<Ԕ�<���<cŃ<`H�<cŃ<���<Ԕ�<A{�<0�<�#�<F��<�R�<T��<�+�<�l�<`   `   '�<���<�U�<�U�<��<�'�<X �<�i�<��<�h�<��z<�Yj<L�d<�Yj<��z<�h�<��<�i�<X �<�'�<��<�U�<�U�<���<`   `   Ni�<��<p2�<��<�u�<#��<�O�<#�<~2�<�&|<�Ha<�dO<TI<�dO<�Ha<�&|<~2�<#�<�O�<#��<�u�<��<p2�<��<`   `   �i�<=
�< ��<���<?�<O��<2A�<z��<�<�Oi<�L<�\9<��2<�\9<�L<�Oi<�<z��<2A�<O��<?�<���< ��<=
�<`   `   �Q�<���<���<�r�<^J�<�>�<f�<���<��<�Y\<��><k�*<��#<k�*<��><�Y\<��<�<f�<�>�<^J�<�r�<���<���<`   `   �F�<���<���<Pd�<�;�<5�<ԁ�<Ï<�Oz<��V<;9<�{%<u�<�{%<;9<��V<�Oz<Ï<ԁ�<5�<�;�<Pd�<���<���<`   `   9s�<�<���<���<K+�<���<Ƒ�<D��<i}{<��Y<t>=<�_*<R�#<�_*<t>=<��Y<h}{<D��<Ƒ�<���<J+�<���<���<�<`   `   ^ �<D��<���<�S�<�;�<c��<���<�<���<�Vd<�aJ<C9<�3<C9<�aJ<�Vd<���<~�<���<c��<�;�<�S�<���<D��<`   `   ��<���<�^�<��<x{�<�5�<��<�"�<终<�v<�X_<�2P<��J<�2P<�X_<�v<终<�"�<��<�5�<x{�<��<�^�<���<`   `   ���<l��<���<u��<eɼ<��<�ĩ<|'�<V�<g��<z<�hm<��h<�hm<z<g��<V�<|'�<�ĩ<��<eɼ<u��<���<l��<`   `   ���<��<���<X��<��<��<Hͯ<���<�ڜ<^��<|�<J	�<�D�<J	�<|�<]��<�ڜ<���<Hͯ<��<��<W��<���<��<`   `   o��<���<]�<L�<���<ν�<ً�<���<�F�<�]�<枛<�͗<w�<�͗<枛<�]�<�F�<���<ً�<ν�<���<L�<\�<���<`   `   d��<mE�<��<���<K5�<���<�}�<���<鎳<;��<坪<&�<���<&�<坪<;��<莳<���<�}�<���<K5�<���<��<mE�<`   `   _
�<��<:T�<n��<��<�h�<���<��<H3�<-@�<P;�<B1�<G-�<B1�<P;�<-@�<G3�<��<���<�h�<��<n��<:T�<��<`   `   ��<=�<��<nz�<�\�<�I�<b.�<
��<U��<#�<�x�<��<���<��<�x�<#�<T��<
��<b.�<�I�<�\�<nz�<��<=�<`   `   ��<�V�<��<�:�<"��<�<�j�<��<��<���<;"�<�{�<&��<�{�<;"�<���<��<��<�j�<�<"��<�:�<��<�V�<`   `   ���<u>�<�=�<8��<��</p�<�K�<A��<qZ�<�l�<�.�<��<��<��<�.�<�l�<qZ�<@��<�K�</p�< ��<8��<�=�<u>�<`   `   (~�<���<Y�<'��<�<@g�<���<���<�q�<���<���<�0�<�a�<�0�<���<���<�q�<���<���<@g�<�<'��<Y�<���<`   `   ��<�6�< ��<���<&�<���<f��<���<%��<x�<>��<� �<R�<� �<>��<x�<%��<���<f��<���<&�<���< ��<�6�<`   `   *��<v�<���< ��<��<j��<z��<�{�<��<���<���<�t�<b��<�t�<���<���<��<�{�<z��<j��<��< ��<���<v�<`   `   ��<+~�<�#�<{��<���<T �<uq�<
w�<Y�<[�<Oe�<Q.�<Pr�<Q.�<Oe�<[�<Y�<
w�<uq�<T �<���<{��<�#�<+~�<`   `   4��<�>�<��<>��<$W�<z	�<���<���<;��<���<�~�<f�<���<f�<�~�<���<;��<���<���<z	�<$W�<>��<��<�>�<`   `   V��<aM�<�c�<)��<�^�<�r�<�h�<���<���<�e�<��<�&�<]��<�&�<��<�e�<���<���<�h�<�r�<�^�<)��<�c�<aM�<`   `   ��<z��<�<��<���<�d�<���<O��<U��<�{�<�\�<���<���<���<�\�<�{�<U��<O��<���<�d�<���<��<�<z��<`   `   ���<��<�:�<�/�<���<���<(��<n��<h�<�2�<=�<���<���<���<=�<�2�<h�<n��<(��<���<���<�/�<�:�<��<`   `   rB�<�G�<�/�<��<Ƽ�<s-�<�U�<���<R��<���<;��<c)�<���<c)�<;��<���<R��<���<�U�<s-�<Ƽ�<��<�/�<�G�<`   `   w�<!(�<KI�<���<���<�[�<z��<��<��<��<��<B}�<���<B}�<��<��<��<��<z��<�[�<���<���<KI�<!(�<`   `   1��<Ӱ�<6��<�ؽ<���<���<�h�<'a�<�v�<���<��<[��<��<[��<��<���<�v�<'a�<�h�<���<���<�ؽ<6��<Ӱ�<`   `   �+�<�U�<���<���<�n�<��<q=�<�9�<�R�<<��<f��<zs�<$��<zs�<f��<<��<�R�<�9�<q=�<��<�n�<���<���<�U�<`   `   �O�<�p�<w��<Tm�<��<d �<8��<[�<�R�<Yr�<���<4C�<���<4C�<���<Yr�<�R�<[�<8��<d �<��<Tm�<w��<�p�<`   `   �%�<l2�</+�<+��<�߿<XT�<�t�<j��<���<F��<���<��<���<��<���<F��<���<j��<�t�<XT�<�߿<+��</+�<l2�<`   `   ���<嗵<W7�<�!�<z��<���<$�<��<QC�<c��<���<��<���<��<���<c��<QC�<��<$�<���<{��<�!�<W7�<嗵<`   `   ���<�k�<���<3޾<W��<t��<7r�<;��<�e�<@��<D�<|]�<a��<|]�<D�<@��<�e�<<��<7r�<t��<W��<3޾<���<�k�<`   `   ��<�Q�<i�<��<���<��<�x�<���<�
�<B��<��<<��<�E�<<��<��<B��<�
�<���<�x�<��<���<��<i�<�Q�<`   `   �j�<���<��<���<h��<D�<}�<���<u/�<`�<aN�<e��<�-�<e��<aN�<`�<u/�<���<}�<D�<h��<���<��<���<`   `   �L�<��<�R�<l�<"��<5��<�<�<	��<'t�<���<Y�<|�<Y�<���<'t�<	��<�<�<5��<"��<l�<�R�<��<`   `   ?��<X�<rw�<���<��<���<_Z�<ݜ�<n��<#��<L��<4�<��<4�<L��<#��<n��<ݜ�<_Z�<���<��<���<rw�<X�<`   `   G-�<B1�<P;�<-@�<G3�<��<���<�h�<��<n��<:T�<��<_
�<��<:T�<n��<��<�h�<���<��<G3�<-@�<P;�<B1�<`   `   ���<��<�x�<#�<T��<
��<a.�<�I�<�\�<nz�<��<=�<��<=�<��<nz�<�\�<�I�<a.�<
��<T��<#�<�x�<��<`   `   &��<�{�<;"�<���<��<��<�j�<�<"��<�:�<��<�V�<��<�V�<��<�:�<"��<�<�j�<��<��<���<;"�<�{�<`   `   ��<��<�.�<�l�<qZ�<@��<�K�</p�< ��<8��<�=�<u>�<���<u>�<�=�<8��< ��</p�<�K�<@��<qZ�<�l�<�.�<��<`   `   �a�<�0�<���<���<�q�<���<���<@g�<�<'��<Y�<���<(~�<���<Y�<'��<�<@g�<���<���<�q�<���<���<�0�<`   `   R�<� �<>��<x�<%��<���<f��<���<&�<���< ��<�6�<��<�6�< ��<���<&�<���<f��<���<%��<x�<>��<� �<`   `   b��<�t�<���<���<��<�{�<z��<j��<��< ��<���<v�<*��<v�<���< ��<��<j��<z��<�{�<��<���<���<�t�<`   `   Pr�<Q.�<Oe�<[�<Y�<
w�<uq�<T �<���<z��<�#�<*~�<��<*~�<�#�<z��<���<S �<tq�<
w�<Y�<[�<Oe�<Q.�<`   `   ���<f�<�~�<���<;��<���<���<z	�<$W�<>��<��<�>�<4��<�>�<��<>��<$W�<z	�<���<���<;��<���<�~�<f�<`   `   ]��<�&�<��<�e�<���<���<�h�<�r�<�^�<)��<�c�<aM�<V��<aM�<�c�<)��<�^�<�r�<�h�<���<���<�e�<��<�&�<`   `   ���<���<�\�<�{�<U��<O��<���<�d�<���<��<�<z��<��<z��<�<��<���<�d�<���<O��<U��<�{�<�\�<���<`   `   ���<���<=�<�2�<h�<n��<(��<���<���<�/�<�:�<��<���<��<�:�<�/�<���<���<(��<n��<h�<�2�<=�<���<`   `   ���<c)�<;��<���<R��<���<�U�<t-�<Ƽ�<��<�/�<�G�<rB�<�G�<�/�<��<Ƽ�<s-�<�U�<���<Q��<���<;��<c)�<`   `   ���<B}�<��<��<��<��<{��<�[�<���<���<KI�<!(�<w�<!(�<KI�<���<���<�[�<z��<��<��<��<��<B}�<`   `   ��<[��<��<���<�v�<(a�<�h�<���<���<�ؽ<6��<Ӱ�<1��<Ӱ�<6��<�ؽ<���<���<�h�<'a�<�v�<���<��<[��<`   `   $��<zs�<f��<=��<�R�<�9�<q=�<��<�n�<���<���<�U�<�+�<�U�<���<���<�n�<��<q=�<�9�<�R�<<��<f��<zs�<`   `   ���<4C�<���<Yr�<�R�<[�<8��<e �<��<Tm�<w��<�p�<�O�<�p�<w��<Tm�<��<d �<8��<[�<�R�<Yr�<���<4C�<`   `   ���<��<���<F��<���<k��<�t�<YT�<�߿<+��</+�<m2�<�%�<l2�</+�<+��<�߿<XT�<�t�<j��<���<F��<���<��<`   `   ���<��<���<c��<RC�<��<$�<���<{��<�!�<W7�<嗵<���<嗵<W7�<�!�<z��<���<$�<��<QC�<c��<���<��<`   `   a��<|]�<D�<@��<�e�<<��<7r�<t��<W��<4޾<���<�k�<���<�k�<���<3޾<W��<t��<7r�<;��<�e�<@��<D�<|]�<`   `   �E�<<��<��<C��<�
�<���<�x�<��<���<��<i�<�Q�<��<�Q�<i�<��<���<��<�x�<���<�
�<B��<��<<��<`   `   �-�<e��<bN�<`�<u/�<���<~�<D�<h��<���<��<���<�j�<���<��<���<h��<D�<}�<���<u/�<`�<aN�<e��<`   `   |�<Y�<���<'t�<
��<�<�<5��<#��<l�<�R�<��<�L�<��<�R�<l�<"��<5��<�<�<	��<'t�<���<Y�<`   `   ��<4�<L��<#��<n��<ݜ�<_Z�<���<��<���<rw�<X�<?��<X�<rw�<���<��<���<_Z�<ݜ�<n��<#��<L��<4�<`   `   ��<��<7��<�w�<=��<���<Xw�<��<��<���<���<q��<C��<q��<���<���<��<��<Xw�<���<=��<�w�<7��<��<`   `    �<�:�<��<��<�	�<�z�<W
�<���<0$�<�u�<9}�<Z%�<	_�<Z%�<9}�<�u�<0$�<���<W
�<�z�<�	�<��<��<�:�<`   `   �j�<מ�<�H�<FT�<���<u/�<���<�c�<���<�,�<�*�<1��<I�<0��<�*�<�,�<���<�c�<���<u/�<���<FT�<�H�<מ�<`   `   ���< 7�<0��<,�<�g�<���<���<�8�<��<5��<��<.u�<5��<.u�<��<4��<��<�8�<���<���<�g�<,�<0��< 7�<`   `   ��<���<ũ�<S��<g6�<���<�y�<~�<�t�<���<d��<��<�@�<��<d��<���<�t�<~�<�y�<���<g6�<S��<ũ�<���<`   `   6��<5��<���<���<��<Ʀ�<G�<���<�)�<�B�<R�<Ԗ�<k��<Ԗ�<R�<�B�<�)�<���<G�<Ʀ�<��<���<���<5��<`   `   ր�<���<�q�<���<���<�r�<��<�|�<���<4��<���<���<�'�<���<���<4��<���<�|�<��<�r�<���<���<�q�<���<`   `   ��<��<o�<�y�<���<�:�<��< �<�:�<�,�<���<�?�<\�<�?�<���<�,�<�:�< �<��<�:�<���<�y�<o�<��<`   `   g��<^��<�m�<�f�<���<���<B�<��<��<Bg�<��<#]�<>u�<#]�<��<Bg�<��<��<B�<���<���<�f�<�m�<^��<`   `   ��<���<�U�<>�<uX�<��<���<U��<^��<�z�<=�<�M�<�f�<�M�<=�<�z�<^��<U��<���<��<uX�<>�<�U�<���<`   `   O�<Z��<��<���<���<���<���<��<z��<�T�<���<P�<��<P�<���<�T�<z��<��<���<���<���<���<��<Z��<`   `   0��<"�<w��<-\�<oD�<0�<�
�<���<mn�<��<�Q�<r��<���<r��<�Q�<��<mn�<���<�
�<0�<oD�<-\�<w��<"�<`   `   �!�<�P�<9��<x��<�\�<%'�<
��<�m�<���<�M�<��<��<p��<��<��<�M�<���<�m�<
��<%'�<�\�<x��<9��<�P�<`   `   �0�<�[�<H��<�|�<�4�<���<.f�<��<#"�<_h�<��<U��<d��<U��<��<_h�<#"�<��<.f�<���<�4�<�|�<H��<�[�<`   `   $�<�?�<Q��<�<�<���<�W�<?��<L��<��<H�<^j�<Y��<s��<Y��<^j�<H�<��<L��<?��<�W�<���<�<�<Q��<�?�<`   `   ���<-�<�m�<���<�S�<���<p��<���<��<���<��<�<-#�<�<��<���<��<���<p��<���<�S�<���<�m�<-�<`   `   -��<F��<�6�<,��<)��<���<i��<��<L��<Y��<�z�<z��<��<z��<�z�<Y��<M��<��<i��<���<)��<,��<�6�<F��<`   `   ���<g��< �<�6�<�<�<��<���<4��<7�<P �<���<��<���<��<���<P �<7�<5��<���<��<�<�<�6�< �<g��<`   `   �-�<(-�<�%�<K
�<���<�k�<W��<�^�<��<w��<�Q�<�>�<�;�<�>�<�Q�<w��<��<�^�<W��<�k�<���<K
�<�%�<(-�<`   `   y��<e��<�Y�<�<���<=��<��<�W�<���<�1�<���<��<���<��<���<�1�<���<�W�<��<=��<���<�<�Y�<e��<`   `   #�<��<:��<\&�<�c�<kx�<�z�<���<x��<��<ը�<Dl�<�[�<Dl�<֨�<��<x��<���<�z�<kx�<�c�<\&�<:��<��<`   `   f��<j��<!'�<lh�<�m�<fJ�<��<���<���<�6�<��<�^�<�E�<�^�<��<�6�<���<���<��<fJ�<�m�<lh�<!'�<j��<`   `   �l�<[;�<3��<-��<T��<�Q�<���<���<Z��<��<S�<S��<M~�<S��<S�<��<Z��<���<���<�Q�<T��<-��<3��<[;�<`   `   ��<���<�=�<�A�<���<��<'�<��<�p�<�l�<��<2�<�	�<2�<��<�l�<�p�<��<'�<��<���<�A�<�=�<���<`   `   C��<q��<���<���<��<��<Xw�<���<=��<�w�<7��<��<��<��<7��<�w�<=��<���<Xw�<��<��<���<���<q��<`   `   	_�<Z%�<9}�<�u�<0$�<���<W
�<�z�<�	�<��<��<�:�< �<�:�<��<��<�	�<�z�<W
�<���<0$�<�u�<9}�<Z%�<`   `   I�<0��<�*�<�,�<���<�c�<���<t/�<���<FT�<�H�<מ�<�j�<מ�<�H�<FT�<���<t/�<���<�c�<���<�,�<�*�<0��<`   `   5��<-u�<��<4��<��<�8�<���<���<�g�<,�<0��< 7�<���< 7�<0��<,�<�g�<���<���<�8�<��<4��<��<-u�<`   `   �@�<��<d��<���<�t�<~�<�y�<���<g6�<S��<ũ�<���<��<���<ũ�<S��<g6�<���<�y�<~�<�t�<���<d��<��<`   `   k��<Ԗ�<R�<�B�<�)�<���<G�<Ʀ�<��<���<���<5��<6��<5��<���<���<��<Ʀ�<G�<���<�)�<�B�<R�<Ԗ�<`   `   �'�<���<���<4��<���<�|�<��<�r�<���<���<�q�<���<ր�<���<�q�<���<���<�r�<��<�|�<���<3��<���<���<`   `   \�<�?�<���<�,�<�:�< �<��<�:�<���<�y�<o�<��<��<��<o�<�y�<���<�:�<��< �<�:�<�,�<���<�?�<`   `   >u�<#]�<��<Bg�<��<��<B�<���<���<�f�<�m�<^��<g��<^��<�m�<�f�<���<���<B�<��<��<Bg�<��<#]�<`   `   �f�<�M�<=�<�z�<^��<U��<���<��<uX�<>�<�U�<���<��<���<�U�<>�<uX�<��<���<T��<^��<�z�<=�<�M�<`   `   ��<P�<���<�T�<z��<��<���<���<���<���<��<Z��<O�<Z��<��<���<���<���<���<��<z��<�T�<���<P�<`   `   ���<r��<�Q�<��<mn�<���<�
�<0�<oD�<-\�<w��<"�<0��<"�<w��<-\�<oD�<0�<�
�<���<mn�<��<�Q�<r��<`   `   q��<��<��<�M�<���<�m�<
��<%'�<�\�<x��<9��<�P�<�!�<�P�<9��<x��<�\�<%'�<
��<�m�<���<�M�<��<��<`   `   d��<U��<��<_h�<$"�<��<.f�<���<�4�<�|�<H��<�[�<�0�<�[�<G��<�|�<�4�<���<.f�<��<#"�<_h�<��<U��<`   `   s��<Y��<^j�<H�<��<L��<?��<�W�<���<�<�<Q��<�?�<$�<�?�<Q��<�<�<���<�W�<?��<L��<��<H�<^j�<Y��<`   `   -#�<�<��<���<��<���<p��<���<�S�<���<�m�<-�<���<-�<�m�<���<�S�<���<p��<���<��<���<��<�<`   `   ��<z��<�z�<Y��<M��<��<i��<���<)��<,��<�6�<F��<-��<F��<�6�<,��<)��<���<i��<��<M��<Y��<�z�<z��<`   `   ���<��<���<Q �<7�<5��<���<��<�<�<�6�< �<g��<���<g��< �<�6�<�<�<��<���<4��<7�<P �<���<��<`   `   �;�<�>�<�Q�<w��<��<�^�<W��<�k�<���<K
�<�%�<)-�<�-�<)-�<�%�<K
�<���<�k�<W��<�^�<��<w��<�Q�<�>�<`   `   ���<��<���<�1�<���<�W�<��<=��<���<�<�Y�<e��<y��<e��<�Y�<�<���<=��<��<�W�<���<�1�<���<��<`   `   �[�<Dl�<֨�<��<x��<���<�z�<kx�<�c�<\&�<:��<��<#�<��<:��<\&�<�c�<kx�<�z�<���<x��<��<֨�<Dl�<`   `   �E�<�^�<��<�6�<���<���<��<fJ�<�m�<mh�<!'�<j��<f��<j��<!'�<lh�<�m�<fJ�<��<���<���<�6�<��<�^�<`   `   M~�<S��<S�<��<Z��<���<���<�Q�<U��<-��<3��<[;�<�l�<[;�<3��<-��<U��<�Q�<���<���<Z��<��<S�<S��<`   `   �	�<2�<��<�l�<�p�<���<'�<��<���<�A�<�=�<���<��<���<�=�<�A�<���<��<'�<��<�p�<�l�<��<2�<`   `   v��<"�<��<��<���<.n�<5�<�<��<~�<���<��<���<��<���<~�<��<�<5�<.n�<���<��<��<"�<`   `   ���<�+�<���<Y��<:��<W�< ��<��<�]�<���<d��<ͼ�<2��<ͼ�<d��<���<�]�<��< ��<W�<:��<Y��<���<�+�<`   `   �n�<��<��<���<��<��<4	�<U��<��<Hg�<�o�<��<BR�<��<�o�<Hg�<��<U��<4	�<��<��<���<��<��<`   `   �2�<^�<Z��< ��<��<z��<�M�<���<N�<r0�<��<���<S��<���<��<r0�<N�<���<�M�<z��<��< ��<Y��<^�<`   `   9H�<"o�<���<:��<��<|��<���<7�<#(�<D+�<Q��<�m�<���<�m�<Q��<D+�<#(�<7�<���<|��<��<:��<���<"o�<`   `   I��<���<1�<���<���<��<ه�<r��<Fx�<�H�<���<�W�<�{�<�W�<���<�H�<Fx�<r��<ه�<��<���<���<1�<���<`   `   �Z�<av�<	��<�C�<l��<���<Xl�<.�<#��<���<�<�\�<y�<�\�<�<���<#��<.�<Xl�<���<l��<�C�<	��<av�<`   `   WM�<=`�<|��<G��<�]�<^��<�i�<���<�q�<��<}1�<?o�<C��<?o�<}1�<��<�q�<���<�i�<^��<�]�<G��<|��<=`�<`   `   �s�<'|�<���<���<{��<`5�<)x�<���<���<4�</b�<���<���<���</b�<4�<���<���<)x�<`5�<{��<���<���<'|�<`   `   z��<���<��<��<���<{��<��<��<�{�<|�<J�<D��<���<D��<J�<|�<�{�<��<��<{��<���<��<��<���<`   `   ��<H��<���<���<N:�<���<���<�,�<)��<��<i�<�f�<Y�<�f�<i�<��<)��<�,�<���<���<N:�<���<���<H��<`   `   �9�<e �<���<W�<r��<�
�<�Y�<$��<"�<l��<�W�<O$�<��<O$�<�W�<l��<"�<$��<�Y�<�
�<r��<W�<���<e �<`   `   F+�<��<m��<���<� �<���<g��<��<�-�<~��<E�</��<���</��<E�<~��<�-�<��<g��<���<� �<���<m��<��<`   `   ���<n��<��<��<���<���<#T�<_�<���<��<�v�<��<���<��<�v�<��<���<_�<#T�<���<���<��<��<n��<`   `   ���<��<��<|��<���<D��<?_�<+��<���<b{�<޵�<t8�<��<t8�<ߵ�<b{�<���<+��<?_�<D��<���<|��<��<��<`   `   ���<�Y�<\��<�U�< ��<���<��<�\�<��<��<���<�6�<E	�<�6�<���<��<��<�\�<��<���< ��<�U�<\��<�Y�<`   `   ���<̉�<N��<�K�<���<���<c��<Y��<���<���<��<{�<l��<{�<��<���<���<Y��<c��<���<���<�K�<N��<̉�<`   `   i��<�G�<YW�<���<��< ��<M��<���<���<�w�<�r�<9��<f��<9��<�r�<�w�<���<���<M��< ��<��<���<YW�<�G�<`   `   y��<���<���<1�<!"�<���<��<���<��<�A�<3�<���<�T�<���<3�<�A�<��<���<��<���<!"�<1�<���<���<`   `   h	�<��<ӫ�<��<��<���<���<d�<$��<=�<���<�P�<��<�P�<���<=�<$��<d�<���<���<��<��<ӫ�<��<`   `   X��<t��<��<|��<��<���<�a�<�C�<sl�<��<X��<;�<���<;�<X��<��<sl�<�C�<�a�<���<��<|��<��<t��<`   `   ��<�9�<9�<���<���<��<�P�<�>�<	r�<���<���<7O�<��<7O�<���<���<	r�<�>�<�P�<��<���<���<9�<�9�<`   `   &<�<���<���<�t�<"��<t��<�e�<�g�<g��<B�<�:�<���<�b�<���<�:�<B�<g��<�g�<�e�<t��<"��<�t�<���<���<`   `   ;��<`��<@��<�a�<ϡ�<i��<���<}��<��<&��<���<�-�<;�<�-�<���<&��<��<}��<���<i��<ϡ�<�a�<@��<`��<`   `   ���<��<���<~�<��<�<5�<.n�<���<��<��<"�<u��<"�<��<��<���<.n�<5�<�<��<~�<���<��<`   `   2��<̼�<d��<���<�]�<��< ��<W�<:��<Y��<���<�+�<���<�+�<���<Y��<:��<W�< ��<��<�]�<���<d��<̼�<`   `   AR�<��<�o�<Hg�<��<U��<4	�<��<��<���<��<��<�n�<��<��<���<��<��<4	�<U��<��<Hg�<�o�<��<`   `   S��<���<��<q0�<M�<���<�M�<z��<��< ��<Y��<^�<�2�<^�<Y��< ��<��<z��<�M�<���<M�<q0�<��<���<`   `   ���<�m�<P��<D+�<#(�<7�<���<|��<��<:��<���<!o�<8H�<!o�<���<:��<��<|��<���<7�<#(�<C+�<P��<�m�<`   `   �{�<�W�<���<�H�<Fx�<r��<ه�<��<���<���<1�<���<I��<���<1�<���<���<��<ه�<r��<Fx�<�H�<���<�W�<`   `   y�<�\�<�<���<#��<.�<Xl�<���<l��<�C�<	��<av�<�Z�<av�<	��<�C�<l��<���<Xl�<.�<#��<���<�<�\�<`   `   C��<?o�<}1�<��<�q�<���<�i�<^��<�]�<G��<|��<=`�<WM�<=`�<|��<G��<�]�<^��<�i�<���<�q�<��<}1�<?o�<`   `   ���<���</b�<4�<���<���<)x�<`5�<{��<���<���<'|�<�s�<'|�<���<���<{��<`5�<)x�<���<���<4�</b�<���<`   `   ���<D��<J�<|�<�{�<��<��<{��<���<��<��<���<z��<���<��<��<���<{��<��<��<�{�<|�<J�<D��<`   `   Y�<�f�<i�<��<)��<�,�<���<���<N:�<���<���<H��<��<H��<���<���<M:�<���<���<�,�<(��<��<i�<�f�<`   `   ��<O$�<�W�<l��<"�<$��<�Y�<�
�<r��<W�<���<e �<�9�<e �<���<W�<r��<�
�<�Y�<$��<"�<l��<�W�<O$�<`   `   ���</��<E�<~��<�-�<��<h��<���<� �<���<m��<��<F+�<��<m��<���<� �<���<g��<��<�-�<~��<E�</��<`   `   ���<��<�v�<��<���<_�<#T�<���<���<��<��<n��<���<n��<��<��<���<���<"T�<_�<���<��<�v�<��<`   `   ��<t8�<ߵ�<b{�<���<+��<?_�<D��<���<|��<��<��<���<��<��<|��<���<D��<?_�<+��<���<b{�<ߵ�<t8�<`   `   F	�<�6�<���<��<��<�\�<��<���< ��<�U�<\��<�Y�<���<�Y�<\��<�U�< ��<���<��<�\�<��<��<���<�6�<`   `   l��<{�<��<���<���<Y��<c��<���<���<�K�<N��<̉�<���<̉�<N��<�K�<���<���<c��<Y��<���<���<��<{�<`   `   f��<9��<�r�<�w�<���<���<M��<��<��<���<YW�<�G�<i��<�G�<YW�<���<��< ��<M��<���<���<�w�<�r�<9��<`   `   �T�<���<3�<�A�<��<���<��<���<""�<1�<���<���<y��<���<���<1�<!"�<���<��<���<��<�A�<3�<���<`   `   ��<�P�<���<=�<$��<d�<���<���<��<��<ӫ�<��<h	�<��<ӫ�<��<��<���<���<d�<$��<=�<���<�P�<`   `   ���<;�<X��<��<tl�<�C�<�a�<���<��<|��<��<t��<X��<t��<��<|��<��<���<�a�<�C�<sl�<��<X��<;�<`   `   ��<7O�<���<���<	r�<�>�<�P�<��<���<���<9�<�9�<��<�9�<9�<���<���<��<�P�<�>�<	r�<���<���<7O�<`   `   �b�<���<�:�<B�<g��<�g�<�e�<t��<"��<�t�<���<���<&<�<���<���<�t�<"��<t��<�e�<�g�<g��<B�<�:�<���<`   `   ;�<�-�<���<&��<��<}��<���<i��<ϡ�<�a�<@��<`��<;��<`��<@��<�a�<ϡ�<i��<���<}��<��<&��<���<�-�<`   `   �
�<�5�<���<W��<��<"�<���<~�<�/�<Ǳ�<O��<���<���<���<O��<Ǳ�<�/�<}�<���<"�<��<W��<���<�5�<`   `   ,�<�S�<���<"��<���<���<oM�<r��<eQ�<V��<{��<�\�<��<�\�<{��<V��<eQ�<r��<oM�<���<���<"��<���<�S�<`   `   d��<K��<�"�<���<Z��<���<'�<�l�<���<���<U��<U�<��<U�<U��<���<���<�l�<'�<���<Z��<���<�"�<K��<`   `   �E�<pd�<���<�X�<�$�<��<A-�<�K�<�_�<OV�<��<f��<C��<f��<��<OV�<�_�<�K�<A-�<��<�$�<�X�<���<pd�<`   `   ,Q�<�j�<˶�<T3�<k��<��<�~�<�k�<%K�<�<��<��<�8�<��<��<�<%K�<�k�<�~�<��<k��<T3�<ʶ�<�j�<`   `   ���<���<� �<�\�<���<=n�<K�<h��<Yp�<�	�<���<���<#��<���<���<�	�<Yp�<h��<K�<=n�<���<�\�<� �<���<`   `   {m�<�x�<ƙ�<��<��<�u�<���<�O�<���<�0�<�<ֽ�<E��<ֽ�<�<�0�<���<�O�<���<�u�<��<��<ƙ�<�x�<`   `   rs�<�u�<�z�<���<���<a��<���<� �<N4�<�i�<���<#��<���<#��<���<�i�<N4�<� �<���<a��<���<���<�z�<�u�<`   `   ���<p��<w��<�l�<{?�<��<���<���<f��<Ŷ�<��<���<(��<���<��<Ŷ�<f��<���<���<��<{?�<�l�<w��<p��<`   `   %�<:�<���<�t�<� �<���<3�<��<�B�<F�<���<���<p��<���<���<F�<�B�<��<3�<���<� �<�t�<���<:�<`   `   9��<�}�<M�<���<���<���<�$�<�d�<��<eD�<,��<!��<˶�<!��<,��<eD�<��<�d�<�$�<���<���<���<M�<�}�<`   `   ��<���<�P�<b}�<9t�<XO�<�'�<��<z&�<k�<���<1��<(��<1��<���<k�<z&�<��<�'�<XO�<9t�<b}�<�P�<���<`   `   u5�<c��<�N�<C�<-��<Sy�<w��<���<>e�<n�<���<�U�<{9�<�U�<���<n�<>e�<���<w��<Sy�<-��<C�<�N�<c��<`   `   J�<L��<���<Ŷ�<n"�<�^�<*��<���<�q�<�D�<�k�<&��<��<&��<�k�<�D�<�q�<���<*��<�^�<n"�<Ŷ�<���<L��<`   `   +o�<��<�/�<���<7��<���<���<���<
E�<���<���<'W�<�+�<'W�<���<���<
E�<���<���<���<7��<���<�/�<��<`   `   *K�<���<��<LS�<�V�<��<6��<Q��<z��<H]�<&F�<k��<h�<k��<&F�<H]�<z��<Q��<6��<��<�V�<LS�<��<���<`   `   {��<�1�<��<g�<G�<���<�|�<�7�<=�<<��<ey�<O��<7��<O��<ey�<<��<=�<�7�<�|�<���<G�<g�<��<�1�<`   `   �H�<��<3��<���<@��<DU�<���<(z�<yl�<���<j��<���<��<���<j��<���<yl�<(z�<���<DU�<@��<���<3��<��<`   `   �x�<��<��<1)�<0��<r�<���<Y��<�y�<���<.��<���<G��<���<.��<���<�y�<Y��<���<r�<0��<1)�<��<��<`   `   �;�<���<_��<���<x��<6S�<8��<���<�u�<g��<d��<L��<���<L��<d��<g��<�u�<���<8��<6S�<x��<���<_��<���<`   `   ��<@S�<�=�<+��<�m�<[�<ê�<�i�<�q�<x��<Ƶ�<��<_��<��<Ƶ�<x��<�q�<�i�<ê�<[�<�m�<+��<�=�<@S�<`   `    ��<���<X��<�<��<���<��<5]�<"��<���<���<XF�<��<XF�<���<���<"��<5]�<��<���<��<�<X��<���<`   `   �1�<I��<���<q�<��<��<�j�<Vn�<˱�<.L�<�J�<ʷ�<��<ʷ�<�J�<.L�<˱�<Vn�<�j�<��<��<q�<���<I��<`   `   �y�<k-�<�P�<d��<�J�<�h�<y|�<���<��<���<���<�X�<>*�<�X�<���<���<��<���<y|�<�h�<�J�<d��<�P�<k-�<`   `   ���<���<O��<Ǳ�<�/�<}�<���<"�<��<W��<���<�5�<�
�<�5�<���<W��<��<"�<���<}�<�/�<Ǳ�<O��<���<`   `   ��<�\�<{��<V��<eQ�<r��<oM�<���<���<"��<���<�S�<,�<�S�<���<"��<���<���<oM�<r��<eQ�<V��<{��<�\�<`   `   ��<U�<U��<���<���<�l�<'�<���<Z��<���<�"�<K��<c��<K��<�"�<���<Z��<���<'�<�l�<���<���<U��<U�<`   `   C��<f��<��<OV�<�_�<�K�<A-�<��<�$�<�X�<���<pd�<�E�<pd�<���<�X�<�$�<��<A-�<�K�<�_�<OV�<��<f��<`   `   �8�<��<��<�<%K�<�k�<�~�<��<k��<T3�<ʶ�<�j�<,Q�<�j�<ʶ�<T3�<k��<��<�~�<�k�<%K�<�<��<��<`   `   #��<���<���<�	�<Yp�<h��<K�<=n�<���<�\�<� �<���<���<���<� �<�\�<���<=n�<K�<h��<Yp�<�	�<���<���<`   `   E��<ֽ�<�<�0�<���<�O�<���<�u�<��<��<ƙ�<�x�<{m�<�x�<ƙ�<��<��<�u�<���<�O�<���<�0�<�<ֽ�<`   `   ���<#��<���<�i�<N4�<� �<���<a��<���<���<�z�<�u�<rs�<�u�<�z�<���<���<a��<���<� �<N4�<�i�<���<#��<`   `   (��<���<��<Ŷ�<f��<���<���<��<{?�<�l�<w��<p��<���<p��<w��<�l�<{?�<��<���<���<f��<Ŷ�<��<���<`   `   p��<���<���<F�<�B�<��<3�<���<� �<�t�<���<:�<%�<:�<���<�t�<� �<���<3�<��<�B�<F�<���<���<`   `   ˶�<!��<,��<eD�<��<�d�<�$�<���<���<���<M�<�}�<9��<�}�<M�<���<���<���<�$�<�d�<��<eD�<,��<!��<`   `   (��<1��<���<k�<z&�<��<�'�<XO�<9t�<b}�<�P�<���<��<���<�P�<b}�<9t�<XO�<�'�<��<z&�<k�<���<1��<`   `   {9�<�U�<���<n�<>e�<���<w��<Sy�<-��<C�<�N�<c��<u5�<c��<�N�<C�<-��<Sy�<v��<���<>e�<n�<���<�U�<`   `   ��<&��<�k�<�D�<�q�<���<*��<�^�<n"�<Ŷ�<���<L��<J�<L��<���<Ŷ�<n"�<�^�<*��<���<�q�<�D�<�k�<&��<`   `   �+�<'W�<���<���<E�<���<���<���<7��<���<�/�<��<+o�<��<�/�<���<7��<���<���<���<
E�<���<���<'W�<`   `   h�<k��<&F�<H]�<z��<R��<6��<��<�V�<MS�<��<���<*K�<���<��<LS�<�V�<��<6��<Q��<z��<H]�<&F�<k��<`   `   7��<O��<ey�<<��<=�<�7�<�|�<���<G�<g�<��<�1�<{��<�1�<��<g�<G�<���<�|�<�7�<=�<<��<ey�<O��<`   `   ��<���<j��<���<zl�<(z�<���<DU�<@��<���<3��<��<�H�<��<3��<���<@��<DU�<���<(z�<yl�<���<j��<���<`   `   G��<���<.��<���<�y�<Y��<���<r�<0��<1)�<��<��<�x�<��<��<1)�<0��<r�<���<Y��<�y�<���<.��<���<`   `   ���<L��<d��<g��<�u�<���<8��<6S�<x��<���<_��<���<�;�<���<_��<���<x��<6S�<8��<���<�u�<g��<d��<L��<`   `   `��<��<Ƶ�<x��<�q�<�i�<ê�<[�<�m�<,��<�=�<@S�<��<@S�<�=�<+��<�m�<[�<ê�<�i�<�q�<x��<Ƶ�<��<`   `   ��<XF�<���<���<"��<5]�<��<���<��<�<X��<���< ��<���<X��<�<��<���<��<5]�<"��<���<���<XF�<`   `   ��<ʷ�<�J�<.L�<˱�<Vn�<�j�<��<��<q�<���<I��<�1�<I��<���<q�<��<��<�j�<Vn�<˱�<.L�<�J�<ʷ�<`   `   >*�<�X�<���<���<��<���<z|�<�h�<�J�<d��<�P�<k-�<�y�<k-�<�P�<d��<�J�<�h�<z|�<���<��<���<���<�X�<`   `   ���<���<��<���<���<���<>�<m��<�
�<�H�<E�<+��<��<+��<E�<�H�<�
�<m��<>�<���<���<���<��<���<`   `   ���<"��<Y+�<f��<$��<S��<���<L�<+4�<�F�<
 �<��<���<��<
 �<�F�<+4�<L�<���<S��<$��<f��<Y+�<"��<`   `   ��<��<�s�<i��<���<���<��<���<���<��<:�<}��<��<}��<:�<��<���<���<��<���<���<i��<�s�<��<`   `   ��<x��<���<�n�<��< ��<��<^r�<�B�<���<Q��<���<!�<���<Q��<���<�B�<^r�<��< ��<��<�n�<���<x��<`   `   �v�<D��<!��<� �<~��<�-�<|��<:�<(�<d��<�3�<;z�<���<;z�<�3�<d��<(�<:�<|��<�-�<~��<� �<!��<D��<`   `    ��<T��<V��<��<{b�<���<dC�<���<�:�<���<~ �<�9�<�L�<�9�<~ �<���<�:�<���<dC�<���<{b�<��<V��<T��<`   `   ��<��<
,�<�E�<dl�<���< ��<�+�<�u�<V��<o��<��<'�<��<o��<V��<�u�<�+�< ��<���<dl�<�E�<
,�<��<`   `   ��<	��<��<���<��<���<���<N��<��<	��<��<��<��<��<��<	��<��<N��<���<���<��<���<��<	��<`   `   _��<��<���<�\�<A�<q��<���<�X�<F:�<�&�<��<��<X�<��<��<�&�<F:�<�X�<���<p��<A�<�\�<���<��<`   `   ��<j��<��<��<���<H�<K��<x
�<ب�<�g�<P:�<N"�<�<N"�<P:�<�g�<ب�<x
�<K��<H�<���<��<��<j��<`   `   ��<���<m��<V��<)�<�R�<�|�<��<��<A��<O�<m �<�<m �<O�<A��<��<��<�|�<�R�<)�<V��<m��<���<`   `   l,�<���<uw�<���<)��<���<^e�<�[�<�x�<���<�R�<'�<���<'�<�R�<���<�x�<�[�<^e�<���<)��<���<uw�<���<`   `   x�<��<�8�<�9�<���<���<R,�<e��<x��<���<]=�<���<���<���<]=�<���<x��<e��<R,�<���<���<�9�<�8�<��<`   `   O��<s�<9��<��<��<pj�<\��<>1�<;��<t��<^�<���<�r�<���<^�<t��<;��<>1�<]��<pj�<��<��<9��<s�<`   `   }��<���<)��<ly�<���<L��<��<IQ�<���<E��<u��<�0�<E�<�0�<u��<E��<���<IQ�<��<L��<���<ly�<)��<���<`   `   ���<b�<�s�<��<�4�<�0�<�#�<c5�<��<B-�<�7�<Z��<�z�<Z��<�7�<B-�<��<c5�<�#�<�0�<�4�<��<�s�<b�<`   `   F��<���<���<#�<�3�<��<���<���<^�<C��<b��<8�<��<8�<b��<C��<^�<���<���<��<�3�<#�<���<���<`   `   ��<Y�<�V�<���<"��<D��<Mg�<�M�<�x�<��<���<�Y�<0%�<�Y�<���<��<�x�<�M�<Mg�<D��<"��<���<�V�<Y�<`   `   ���<���<O��<�<S�<n��<���<���<B��<`D�<�6�<k��<rg�<k��<�6�<`D�<B��<���<���<n��<S�<�<O��<���<`   `   ��<���<Q��<� �<��<���<���<h��<1��<�}�<|w�<���<���<���<|w�<�}�<1��<h��<���<���<��<� �<Q��<���<`   `   	o�<o�<[,�<6��<���<���<���<~��<]�<���<+��<�0�<���<�0�<+��<���<]�<~��<���<���<���<6��<[,�<o�<`   `   ���<���<���<�N�<���<U��<��<���<LO�<��<L#�</��<i�</��<L#�<��<LO�<���<��<U��<���<�N�<���<���<`   `   �1�<��<��<���<cL�<��<��<�<o��<s�<*��<��<d��<��<*��<s�<o��<�<��<��<cL�<���<��<��<`   `   ���<�V�<1��<X��<��<f��<���<sg�<Q�<�<ZH�<��<���<��<ZH�<�<Q�<sg�<���<f��<��<X��<1��<�V�<`   `   ��<+��<E�<�H�<�
�<m��<>�<���<���<���<��<���<���<���<��<���<���<���<>�<m��<�
�<�H�<E�<+��<`   `   ���<��<
 �<�F�<+4�<L�<���<S��<$��<f��<Y+�<"��<���<"��<Y+�<f��<$��<S��<���<L�<+4�<�F�<
 �<��<`   `   ��<}��<:�<��<���<���<��<���<���<i��<�s�<��<��<��<�s�<i��<���<���<��<���<���<��<:�<}��<`   `   !�<���<Q��<���<�B�<^r�<��< ��<��<�n�<���<x��<��<x��<���<�n�<��< ��<��<^r�<�B�<���<Q��<���<`   `   ���<;z�<�3�<d��<(�<:�<|��<�-�<~��<� �<!��<C��<�v�<C��<!��<� �<~��<�-�<|��<:�<(�<d��<�3�<;z�<`   `   �L�<�9�<~ �<���<�:�<���<dC�<���<{b�<��<V��<T��< ��<T��<V��<��<{b�<���<dC�<���<�:�<���<~ �<�9�<`   `   '�<��<o��<V��<�u�<�+�< ��<���<dl�<�E�<
,�<��<��<��<
,�<�E�<dl�<���< ��<�+�<�u�<V��<o��<��<`   `   ��<��<��<	��<��<N��<���<���<��<���<��<	��<��<	��<��<���<��<���<���<N��<��<	��<��<��<`   `   X�<��<��<�&�<F:�<�X�<���<p��<A�<�\�<���<��<^��<��<���<�\�<A�<p��<���<�X�<F:�<�&�<��<��<`   `   �<N"�<P:�<�g�<ب�<x
�<K��<H�<���<��<��<j��<��<j��<��<��<���<H�<K��<x
�<ب�<�g�<P:�<N"�<`   `   �<m �<O�<A��<��<��<�|�<�R�<)�<V��<m��<���<��<���<m��<V��<)�<�R�<�|�<��<��<A��<O�<m �<`   `   ���<'�<�R�<���<�x�<�[�<^e�<���<)��<���<uw�<���<l,�<���<uw�<���<)��<���<^e�<�[�<�x�<���<�R�<'�<`   `   ���<���<]=�<���<x��<e��<R,�<���<���<�9�<�8�<��<x�<��<�8�<�9�<���<���<R,�<e��<x��<���<]=�<���<`   `   �r�<���<^�<u��<;��<>1�<]��<pj�<��<��<9��<s�<O��<s�<9��<��<��<pj�<\��<>1�<;��<t��<^�<���<`   `   E�<�0�<u��<E��<���<IQ�<��<L��<���<ly�<)��<���<}��<���<)��<ly�<���<L��<��<IQ�<���<E��<u��<�0�<`   `   �z�<Z��<�7�<B-�<��<c5�<�#�<�0�<�4�<��<�s�<b�<���<b�<�s�<��<�4�<�0�<�#�<c5�<��<B-�<�7�<Z��<`   `   ��<8�<c��<D��<^�<���<���<��<�3�<#�<���<���<F��<���<���<#�<�3�<��<���<���<^�<C��<c��<8�<`   `   0%�<�Y�<���<��<�x�<�M�<Mg�<E��<"��<���<�V�<Y�<��<Y�<�V�<���<"��<D��<Mg�<�M�<�x�<��<���<�Y�<`   `   rg�<k��<�6�<`D�<B��<���<���<n��<S�<�<O��<���<���<���<O��<�<S�<n��<���<���<B��<`D�<�6�<k��<`   `   ���<���<|w�<�}�<1��<h��<���<���<��<� �<Q��<���<��<���<Q��<� �<��<���<���<h��<1��<�}�<|w�<���<`   `   ���<�0�<+��<���<]�<~��<���<���<���<6��<[,�<o�<	o�<o�<[,�<6��<���<���<���<~��<]�<���<+��<�0�<`   `   i�</��<L#�<��<LO�<���<��<U��<���<�N�<���<���<���<���<���<�N�<���<U��<��<���<LO�<��<L#�</��<`   `   d��<��<*��<s�<o��<�<��<��<cL�<���<��<��<�1�<��<��<���<cL�<��<��<�<o��<s�<*��<��<`   `   ���<��<ZH�<�<Q�<sg�<���<f��<��<Y��<2��<�V�<���<�V�<1��<Y��<��<f��<���<sg�<Q�<�<ZH�<��<`   `   ��<��<��<܈�<3H�<�2�<q;�<�K�<�\�<�O�<.�<��<Z��<��<.�<�O�<�\�<�K�<q;�<�2�<3H�<܈�<��<��<`   `   ���<ո�<��<M��<1)�<���<��<S��<��<���<�%�<H��<���<H��<�%�<���<��<S��<��<���<1)�<M��<��<ո�<`   `   y��<%��<�=�<k��<\8�<���<<��<�s�<�8�<*��<�q�<��<���<��<�q�<*��<�8�<�s�<<��<���<\8�<k��<�=�<%��<`   `   ca�<t�<��<��<	x�<��<��<rK�<���<z�<���<33�<�K�<33�<���<z�<���<qK�<��<��<	x�<��<��<t�<`   `   c�<	#�<�K�<w��<��<;V�<Z��<�P�<���<�;�<���<���<���<���<���<�;�<���<�P�<Z��<;V�<��<w��<�K�<	#�<`   `   �<P
�<�#�<�N�<ˉ�<���<�%�<�~�<%��<�%�<�d�<��<?��<��<�d�<�%�<%��<�~�<�%�<���<ˉ�<�N�<�#�<P
�<`   `   Y%�<t*�<�2�<�A�<bX�<�x�<��<���<m �<�/�<uU�<^n�<Hx�<^n�<uU�<�/�<m �<���<��<�x�<bX�<�A�<�2�<t*�<`   `   �}�<5y�<�m�<�\�<�P�<�C�<�;�<><�<XD�<�P�<%\�<ze�<�i�<ze�<%\�<�P�<XD�<><�<�;�<�C�<�P�<�\�<�m�<5y�<`   `   ��<?��<���<]��<	e�<�$�<���<��<ۘ�<��<�p�<�i�<Gg�<�i�<�p�<��<ۘ�<��<���<�$�<	e�<]��<���<?��<`   `   ���<��<�\�<��<I��<w�<��<HH�<K��<x��<���<bq�<wh�<bq�<���<x��<K��<HH�<��<w�<I��<��<�\�<��<`   `   6^�<wA�<`��<nk�<e��<?�<Pl�<���<kM�<���<���<�r�<�c�<�r�<���<���<kM�<���<Pl�<?�<e��<nk�<`��<wA�<`   `   �<���<�r�<���<��<��<7#�<L�<���<F�<��<�h�<�T�<�h�<��<F�<���<L�<7#�<��<��<���<�r�<���<`   `   ��<�Z�<*��<��<��<���<���<���<h��<��<ؚ�<�M�<14�<�M�<ؚ�<��<h��<���<���<���<��<��<*��<�Z�<`   `   ���<`��<r��<��<��<���<F9�<���<���<��<�x�<��<.��<��<�x�<��<���<���<F9�<���<��<��<r��<`��<`   `   ���<;��<���<6��<{�<4 �<R��<p�<���<���<�=�<w��<c��<w��<�=�<���<���<p�<R��<4 �<{�<6��<���<;��<`   `   �b�<�!�<�d�<�?�<���<�2�<!��<�	�<��<���<x��<_s�<�L�<_s�<x��<���<��<�	�<!��<�2�<���<�?�<�d�<�!�<`   `   <��<IQ�<q��<(V�<Q��<V �<�g�<���<�c�<�I�<�z�<��<���<��<�z�<�I�<�c�<���<�g�<V �<Q��<(V�<q��<IQ�<`   `   �a�<��<bP�<��<��<o��<D�<a�<|��<��<%��<�y�<�N�<�y�<%��<��<|��<a�<D�<o��<��<��<bP�<��<`   `   ��<���<f��<=��<H��<;�<By�<���<c�<T@�<k�<���<���<���<k�<T@�<c�<���<By�<;�<H��<=��<f��<���<`   `   ��<(��<a��<���<*�<�|�<���<�*�<��<b��<#��<zZ�<v0�<zZ�<#��<b��<��<�*�<���<�|�<*�<���<a��<(��<`   `   ~��<W��<=��<Ш�<�8�<��<���<�v�<�&�<��<�J�<#��<=��<#��<�J�<��<�&�<�v�<���<��<�8�<Ш�<=��<W��<`   `   ���<4E�<,��<��<�1�<r��<�0�<���<��<��<c��<}Z�<�4�<}Z�<c��<��<��<���<�0�<r��<�1�<��<,��<4E�<`   `   C.�<C��<�X�<fa�<�)�<���<&m�<�$�<���<��<�d�<���<��<���<�d�<��<���<�$�<&m�<���<�)�<fa�<�X�<C��<`   `   ���<V��<x%�<�H�<N3�<[��<���<��<Ց�<��<=�<��<y��<��<=�<��<Ց�<��<���<[��<N3�<�H�<x%�<V��<`   `   Z��<��<.�<�O�<�\�<�K�<q;�<�2�<2H�<܈�<��<��<��<��<��<܈�<2H�<�2�<q;�<�K�<�\�<�O�<.�<��<`   `   ���<H��<�%�<���<��<S��<��<���<0)�<M��<��<ո�<���<ո�<��<M��<0)�<���<��<S��<��<���<�%�<H��<`   `   ���<��<�q�<*��<�8�<�s�<<��<���<\8�<k��<�=�<%��<y��<%��<�=�<k��<\8�<���<<��<�s�<�8�<*��<�q�<��<`   `   �K�<33�<���<z�<���<qK�<��<��<	x�<��<��<t�<ca�<t�<��<��<	x�<��<��<qK�<���<z�<���<33�<`   `   ���<���<���<�;�<���<�P�<Z��<;V�<��<w��<�K�<	#�<c�<	#�<�K�<w��<��<;V�<Z��<�P�<���<�;�<���<���<`   `   ?��<��<�d�<�%�<%��<�~�<�%�<���<ˉ�<�N�<�#�<P
�<�<P
�<�#�<�N�<ˉ�<���<�%�<�~�<%��<�%�<�d�<��<`   `   Hx�<^n�<uU�<�/�<m �<���<��<�x�<bX�<�A�<�2�<t*�<Y%�<t*�<�2�<�A�<bX�<�x�<��<���<m �<�/�<uU�<^n�<`   `   �i�<ze�<%\�<�P�<XD�<><�<�;�<�C�<�P�<�\�<�m�<5y�<�}�<5y�<�m�<�\�<�P�<�C�<�;�<><�<XD�<�P�<%\�<ze�<`   `   Gg�<�i�<�p�<��<ۘ�<��<���<�$�<	e�<]��<���<?��<��<?��<���<]��<	e�<�$�<���<��<ۘ�<��<�p�<�i�<`   `   wh�<bq�<���<x��<K��<HH�<��<w�<I��<��<�\�<��<���<��<�\�<��<I��<w�<��<HH�<K��<x��<���<bq�<`   `   �c�<�r�<���<���<kM�<���<Pl�<?�<e��<nk�<`��<wA�<6^�<wA�<`��<nk�<e��<?�<Pl�<���<kM�<���<���<�r�<`   `   �T�<�h�<��<F�<���<L�<7#�<��<��<���<�r�<���<�<���<�r�<���<��<��<7#�<L�<���<F�<��<�h�<`   `   14�<�M�<ؚ�<��<h��<���<���<���<��<��<*��<�Z�<��<�Z�<*��<��<��<���<���<���<h��<��<ؚ�<�M�<`   `   .��<��<�x�<��<���<���<F9�<���<��<��<r��<`��<���<`��<r��<��<��<���<F9�<���<���<��<�x�<��<`   `   c��<w��<�=�<���<���<p�<R��<4 �<{�<6��<���<;��<���<;��<���<6��<{�<4 �<R��<p�<���<���<�=�<w��<`   `   �L�<_s�<x��<���<��<�	�<!��<�2�<���<�?�<�d�<�!�<�b�<�!�<�d�<�?�<���<�2�<!��<�	�<��<���<x��<_s�<`   `   ���<��<�z�<�I�<�c�<���<�g�<V �<Q��<(V�<q��<JQ�<<��<IQ�<q��<(V�<Q��<V �<�g�<���<�c�<�I�<�z�<��<`   `   �N�<�y�<%��<��<}��<a�<D�<o��<��<��<bP�<��<�a�<��<bP�<��<��<o��<D�<a�<|��<��<%��<�y�<`   `   ���<���<k�<T@�<c�<���<By�<;�<H��<=��<f��<���<��<���<f��<=��<H��<;�<By�<���<c�<T@�<k�<���<`   `   v0�<zZ�<#��<b��<��<�*�<���<�|�<*�<���<a��<(��<��<(��<a��<���<*�<�|�<���<�*�<��<b��<#��<zZ�<`   `   =��<#��<�J�<��<�&�<�v�<���<��<�8�<Ш�<=��<W��<~��<W��<=��<Ш�<�8�<��<���<�v�<�&�<��<�J�<#��<`   `   �4�<}Z�<c��<��<��<���<�0�<r��<�1�<��<,��<4E�<���<4E�<,��<��<�1�<r��<�0�<���<��<��<c��<}Z�<`   `   ��<���<�d�<��<���<�$�<&m�<���<�)�<fa�<�X�<C��<C.�<C��<�X�<fa�<�)�<���<&m�<�$�<���<��<�d�<���<`   `   y��<��<=�<��<Ց�<��<���<[��<N3�<�H�<x%�<V��<���<V��<x%�<�H�<N3�<[��<���<��<Ց�<��<=�<��<`   `   ��<U#�<h�<0��<Wl�<�!�<���<��<���<�?�<���<g*�<QI�<g*�<���<�?�<���<��<���<�!�<Wl�<0��<h�<U#�<`   `   �<�2�<�n�<��<�R�<���<���<>V�<��<_��<c�<Kl�<��<Kl�<c�<_��<��<>V�<���<���<�R�<��<�n�<�2�<`   `   @W�<�h�<���<S��<�]�<i��<�v�<��<ɤ�<�'�<׎�<���<Z��<���<׎�<�'�<ɤ�<��<�v�<i��<�]�<S��<���<�h�<`   `   F��<z��<y��<�3�<���<���<jq�<:��<[f�<b��<�$�<Z�<�l�<Z�<�$�<b��<Zf�<:��<jq�<���<���<�3�<y��<z��<`   `   LF�<�P�<�n�<۠�< ��<�4�<���<���<DK�<K��<g��<��<W�<��<g��<K��<DK�<���<���<�4�< ��<۠�<�n�<�P�<`   `   `��<��<�< 6�<I`�<���<���<��<O�<���<޴�<���<k��<���<޴�<���<O�<��<���<���<I`�< 6�<�<��<`   `   ���<���<��<��<��<�<�-�<FM�<Dm�<��< ��<7��<]��<7��< ��<��<Dm�<FM�<�-�<�<��<��<��<���<`   `   ���<���<���<d��<��<$��<Ϥ�<���<ɠ�<
��<���<H��<+��<H��<���<
��<ɠ�<���<Ϥ�<$��<��<d��<���<���<`   `   ��<P�<e��<���<��<�]�<-�<�<P��<��<m��<���<��<���<m��<��<P��<�<-�<�]�<��<���<e��<P�<`   `   �C�<b8�<��<f��<Ct�<��<��<(m�<�'�<���<��<���<g��<���<��<���<�'�<(m�<��<��<Ct�<f��<��<b8�<`   `   ���<om�<<.�<R��<�Z�<<��<,R�<s��<�m�<1�<���<b��<��<b��<���<1�<�m�<s��<,R�<<��<�Z�<R��<<.�<om�<`   `   6��<#��<�L�<#��<B2�<V��<W��<I8�<d��<�8�<���<���<���<���<���<�8�<d��<I8�<W��<V��<B2�<#��<�L�<#��<`   `   ���<���<R�<ݸ�<���<�%�< Q�<���<v��<�I�<���<���<z��<���<���<�I�<v��<���< Q�<�%�<���<ݸ�<R�<���<`   `   ��<ڠ�<b-�<F{�<X��<+��<.��<'��<���<*G�<~��<j��<!j�<j��<~��<*G�<���<'��<.��<+��<X��<F{�<b-�<ڠ�<`   `   [�<"S�<g��<�
�<^�<���<z��<���<O��<�-�<���<P�<P4�<P�<���<�-�<O��<���<z��<���<^�<�
�<g��<"S�<`   `   ���<
��<�5�<�\�<aL�<��<m��<��<���<,��<�e�<Q
�<x��<Q
�<�e�<,��<���<��<m��<��<aL�<�\�<�5�<
��<`   `   ��<���<Q�<xm�<O�<m�<��<	��<a��<U��<M�<��<���<��<M�<U��<a��<	��<��<m�<O�<xm�<Q�<���<`   `   ���<���<S&�<�=�<��<A��<ن�<�O�<v:�<?Y�<д�<]P�</�<]P�<д�<?Y�<v:�<�O�<ن�<A��<��<�=�<S&�<���<`   `   ͂�<(O�<��<���<H��<�h�<�!�<b��<���<`��<'J�<I��<���<I��<'J�<`��<���<b��<�!�<�h�<H��<���<��<(O�<`   `   i��<��<��<�5�<��<K��<`��<�i�<TZ�<`}�<���<x�<mW�<x�<���<`}�<TZ�<�i�<`��<K��<��<�5�<��<��<`   `   	�<:��<]K�<�t�<�f�<;�<e�<���<���<U
�<n�<:�<���<:�<n�<U
�<���<���<e�<;�<�f�<�t�<]K�<:��<`   `   �<���<�g�<���<��<���<-n�<[�<g�<���<��<���<��<���<��<���<g�<[�<-n�<���<��<���<�g�<���<`   `   U�<,��<4|�<���<���<��<��<G��<���<ZD�<Ի�<vh�<L�<vh�<Ի�<ZD�<���<G��<��<��<���<���<4|�<,��<`   `   �%�<R�<���<)��<?-�<�D�<�V�<�r�<���<���<Ԃ�<�6�<��<�6�<Ԃ�<���<���<�r�<�V�<�D�<?-�<)��<���<R�<`   `   QI�<g*�<���<�?�<���<��<���<�!�<Wl�</��<h�<U#�<��<U#�<h�</��<Wl�<�!�<���<��<���<�?�<���<g*�<`   `   ��<Kl�<c�<_��<��<>V�<���<���<�R�<��<�n�<�2�<�<�2�<�n�<��<�R�<���<���<>V�<��<_��<c�<Kl�<`   `   Z��<���<׎�<�'�<ɤ�<��<�v�<i��<�]�<S��<���<�h�<@W�<�h�<���<S��<�]�<i��<�v�<��<ɤ�<�'�<׎�<���<`   `   �l�<Z�<�$�<b��<Zf�<:��<jq�<���<���<�3�<y��<z��<F��<z��<y��<�3�<���<���<jq�<:��<Zf�<b��<�$�<Z�<`   `   W�<��<g��<K��<DK�<���<���<�4�< ��<۠�<�n�<�P�<LF�<�P�<�n�<۠�< ��<�4�<���<���<DK�<K��<g��<��<`   `   k��<���<޴�<���<O�<��<���<���<I`�< 6�<�<��<`��<��<�< 6�<I`�<���<���<��<O�<���<޴�<���<`   `   ]��<7��< ��<��<Dm�<FM�<�-�<�<��<��<��<���<���<���<��<��<��<�<�-�<FM�<Dm�<��< ��<7��<`   `   +��<H��<���<
��<ɠ�<���<Ϥ�<$��<��<d��<���<���<���<���<���<d��<��<$��<Ϥ�<���<ɠ�<
��<���<H��<`   `   ��<���<m��<��<P��<�<-�<�]�<��<���<e��<P�<��<P�<e��<���<��<�]�<-�<�<P��<��<m��<���<`   `   g��<���<��<���<�'�<(m�<��<��<Ct�<f��<��<b8�<�C�<b8�<��<f��<Ct�<��<��<(m�<�'�<���<��<���<`   `   ��<b��<���<1�<�m�<s��<,R�<<��<�Z�<R��<<.�<om�<���<om�<<.�<R��<�Z�<<��<,R�<s��<�m�<1�<���<b��<`   `   ���<���<���<�8�<d��<I8�<W��<V��<B2�<$��<�L�<#��<6��<#��<�L�<#��<B2�<V��<W��<I8�<d��<�8�<���<���<`   `   z��<���<���<�I�<v��<���< Q�<�%�<���<ݸ�<R�<���<���<���<R�<ݸ�<���<�%�< Q�<���<v��<�I�<���<���<`   `   !j�<j��<~��<*G�<���<'��<.��<+��<X��<F{�<b-�<ڠ�<��<ڠ�<b-�<F{�<X��<+��<.��<'��<���<*G�<~��<j��<`   `   P4�<P�<���<�-�<O��<���<z��<���<^�<�
�<g��<"S�<[�<"S�<g��<�
�<^�<���<z��<���<O��<�-�<���<P�<`   `   y��<Q
�<�e�<,��<���<��<m��<��<aL�<�\�<�5�<
��<���<
��<�5�<�\�<aL�<��<m��<��<���<,��<�e�<Q
�<`   `   ���<��<M�<U��<a��<	��<��<m�<O�<xm�<Q�<���<��<���<Q�<xm�<O�<m�<��<	��<a��<U��<M�<��<`   `   /�<]P�<д�<?Y�<v:�<�O�<ن�<A��<��<�=�<S&�<���<���<���<S&�<�=�<��<A��<ن�<�O�<v:�<?Y�<д�<]P�<`   `   ���<I��<(J�<`��<���<b��<�!�<�h�<H��<���<��<(O�<͂�<(O�<��<���<H��<�h�<�!�<b��<���<`��<(J�<I��<`   `   mW�<x�<���<`}�<TZ�<�i�<`��<K��<��<�5�<��<��<i��<��<��<�5�<��<K��<`��<�i�<TZ�<`}�<���<x�<`   `   ���<:�<n�<U
�<���<���<e�<;�<�f�<�t�<]K�<:��<
�<:��<]K�<�t�<�f�<;�<e�<���<���<U
�<n�<:�<`   `   ��<���<��<���<g�<[�<-n�<���<��<���<�g�<���<�<���<�g�<���<��<���<-n�<[�<g�<���<��<���<`   `   L�<vh�<Ի�<ZD�<���<G��<��<��<���<���<4|�<,��<U�<,��<4|�<���<���<��<��<G��<���<ZD�<Ի�<vh�<`   `   ��<�6�<Ԃ�<���<���<�r�<�V�<�D�<@-�<)��<���<R�<�%�<R�<���<)��<@-�<�D�<�V�<�r�<���<���<Ԃ�<�6�<`   `   �5�<�G�<�|�<��<�F�<!��<�j�<�	�<���<�(�<N��<���<x��<���<N��<�(�<���<�	�<�j�<!��<�F�<��<�|�<�G�<`   `   RD�< S�<���<G��<2�<#��<�/�<���<�<�<ұ�<��<"G�<^[�<"G�<��<ұ�<�<�<���<�/�<#��<2�<G��<���< S�<`   `   �p�<}�<u��<(��<�8�<j��<��<��<���<�S�<@��<E��<|��<E��<@��<�S�<���<��<��<j��<�8�<(��<u��<}�<`   `   3��<���<���<��<]�<���<=
�<*g�<���<�<�M�<�u�<��<�u�<�M�<�<���<*g�<=
�<���<]�<��<���<���<`   `   �(�<<1�<�H�<�m�<���<���<8 �<me�<���<��<��<�3�<�=�<�3�<��<��<���<me�<8 �<���<���<�m�<�H�<<1�<`   `    ��<	��<���<���<���<%�<�O�<)}�<o��<���<���<	�<"�<	�<���<���<o��<)}�<�O�<%�<���<���<���<	��<`   `   �b�<d�<5g�<'n�<�w�<���<��<Y��<X��<D��<v��<���<O��<���<v��<D��<X��<Y��<��<���<�w�<'n�<5g�<d�<`   `   v)�<�&�<��<�<��<]��<���<6��<���<k��<��<��<e��<��<��<k��<���<6��<���<]��<��<�<��<�&�<`   `   ��<���<���<���<���<�~�<�W�<�4�<��<"�< ��<���<:��<���< ��<"�<��<�4�<�W�<�~�<���<���<���<���<`   `   ���<d��<��<$��<�O�<�<���<ą�<mN�<b"�<|�<���<��<���<|�<b"�<mN�<ą�<���<�<�O�<$��<��<d��<`   `   B��<G��<���<_R�<���<ݗ�<�3�<J��<��<�A�<�<
��<���<
��<�<�A�<��<J��<�3�<ݗ�<���<_R�<���<G��<`   `   ���<-��<i�<0�<Л�<��<u��<��<n��<�Z�<4�<���<���<���<4�<�Z�<n��<��<u��<��<Л�<0�<i�<-��<`   `   3��<�k�<�%�<@��<),�<1��<7��<�[�<���<�i�<��<���<���<���<��<�i�<���<�[�<7��<1��<),�<@��<�%�<�k�<`   `   �0�<��<���<C�<���<���<5�<
��<���<�i�<D�<8��<��<8��<D�<�i�<���<
��<5�<���<���<C�<���<��<`   `   +��<s��<�7�<$��<P��<h+�<�\�<V��<��<�X�<H��<g��<l��<g��<H��<�X�<��<V��<�\�<h+�<P��<$��<�7�<s��<`   `   J�<R��<W~�<7��<p!�<mF�<�e�<��<���<.5�<���<�z�<gb�<�z�<���<.5�<���<��<�e�<mF�<p!�<7��<W~�<R��<`   `   1�<���<]��<q��<�#�<E=�<yP�<�n�<å�<X �<���<�;�<�"�<�;�<���<X �<å�<�n�<yP�<E=�<�#�<q��<]��<���<`   `   /�<���<�s�<���<���<��<�<E5�<#g�<!��<�>�<���<��<���<�>�<!��<#g�<E5�<�<��<���<���<�s�<���<`   `   T��<��<p&�<؀�<��<���<	��<m��<N�<�m�<`��<���<���<���<`��<�m�<N�<m��<	��<���<��<؀�<p&�<��<`   `    =�<��<��<u�<�C�<\�<nn�<Պ�<̾�<�<{��<�M�<�3�<�M�<{��<�<̾�<Պ�<nn�<\�<�C�<u�<��<��<`   `   ���<?��<� �<���<���<���<* �<�%�<�a�<\��<(H�<��<���<��<(H�<\��<�a�<�%�<+ �<���<���<���<� �<?��<`   `   ���<���<w|�<���<�3�<�d�<w��<J��<��<en�<J��<���<���<���<J��<en�<��<J��<w��<�d�<�3�<���<w|�<���<`   `   �C�<�&�<���<�L�<��<;��<�<�`�<��<t'�<ǽ�<}�<{f�<}�<ǽ�<t'�<��<�`�<�<;��<��<�L�<���<�&�<`   `   Α�<�w�<R+�<ų�<@�<o�<���<S�<?t�<K��<B��<�V�<@B�<�V�<B��<K��<?t�<S�<���<o�<@�<ų�<R+�<�w�<`   `   x��<���<N��<�(�<���<�	�<�j�<!��<�F�<��<�|�<�G�<�5�<�G�<�|�<��<�F�<!��<�j�<�	�<���<�(�<N��<���<`   `   ^[�<"G�<��<ұ�<�<�<���<�/�<#��<2�<G��<���< S�<RD�< S�<���<G��<2�<#��<�/�<���<�<�<ұ�<��<"G�<`   `   |��<E��<@��<�S�<���<��<��<j��<�8�<(��<u��<}�<�p�<}�<u��<(��<�8�<j��<��<��<���<�S�<@��<E��<`   `   ��<�u�<�M�<�<���<*g�<=
�<���<]�<��<���<���<3��<���<���<��<]�<���<=
�<*g�<���<�<�M�<�u�<`   `   �=�<�3�<��<��<���<me�<8 �<���<���<�m�<�H�<<1�<�(�<<1�<�H�<�m�<���<���<8 �<me�<���<��<��<�3�<`   `   "�<	�<���<���<o��<)}�<�O�<%�<���<���<���<	��< ��<	��<���<���<���<%�<�O�<)}�<o��<���<���<	�<`   `   O��<���<v��<D��<X��<Y��<��<���<�w�<'n�<5g�<d�<�b�<d�<5g�<'n�<�w�<���<��<Y��<X��<D��<v��<���<`   `   e��<��<��<k��<���<6��<���<]��<��<�<��<�&�<v)�<�&�<��<�<��<]��<���<6��<���<k��<��<��<`   `   :��<���< ��<"�<��<�4�<�W�<�~�<���<���<���<���<��<���<���<���<���<�~�<�W�<�4�<��<"�< ��<���<`   `   ��<���<|�<b"�<mN�<ą�<���<�<�O�<$��<��<d��<���<d��<��<$��<�O�<�<���<ą�<mN�<b"�<|�<���<`   `   ���<
��<�<�A�<��<J��<�3�<ݗ�<���<_R�<���<G��<B��<G��<���<_R�<���<ݗ�<�3�<J��<��<�A�<�<
��<`   `   ���<���<4�<�Z�<n��<��<u��<��<Л�<0�<i�<-��<���<-��<i�<0�<Л�<��<u��<��<n��<�Z�<4�<���<`   `   ���<���<��<�i�<���<�[�<7��<1��<),�<@��<�%�<�k�<3��<�k�<�%�<@��<),�<1��<7��<�[�<���<�i�<��<���<`   `   ��<8��<D�<�i�<���<
��<5�<���<���<C�<���<��<�0�<��<���<C�<���<���<5�<
��<���<�i�<D�<8��<`   `   l��<g��<H��<�X�<��<V��<�\�<h+�<P��<$��<�7�<s��<+��<s��<�7�<$��<P��<h+�<�\�<V��<��<�X�<H��<g��<`   `   gb�<�z�<���</5�<���<��<�e�<mF�<p!�<7��<W~�<R��<J�<R��<W~�<7��<p!�<mF�<�e�<��<���<.5�<���<�z�<`   `   �"�<�;�<���<X �<å�<�n�<yP�<E=�<�#�<q��<]��<���<1�<���<]��<q��<�#�<E=�<yP�<�n�<å�<X �<���<�;�<`   `   ��<���<�>�<!��<#g�<E5�<�<��<���<���<�s�<���</�<���<�s�<���<���<��<�<E5�<#g�<!��<�>�<���<`   `   ���<���<a��<�m�<N�<m��<	��<���<��<؀�<p&�<��<T��<��<p&�<؀�<��<���<	��<m��<N�<�m�<`��<���<`   `   �3�<�M�<{��<�<̾�<Պ�<nn�<\�<�C�<u�<��<��< =�<��<��<u�<�C�<\�<nn�<Պ�<̾�<�<{��<�M�<`   `   ���<��<(H�<\��<�a�<�%�<+ �<���<���<���<� �<?��<���<?��<� �<���<���<���<+ �<�%�<�a�<\��<(H�<��<`   `   ���<���<J��<en�<��<J��<w��<�d�<�3�<���<w|�<���<���<���<w|�<���<�3�<�d�<w��<J��<��<en�<J��<���<`   `   |f�<}�<Ƚ�<t'�<��<�`�<�<;��<��<�L�<���<�&�<�C�<�&�<���<�L�<��<;��<�<�`�<��<t'�<Ƚ�<}�<`   `   @B�<�V�<B��<K��<?t�<S�<���<o�<@�<ų�<S+�<�w�<Α�<�w�<S+�<ų�<@�<o�<���<S�<?t�<K��<B��<�V�<`   `   ��<C$�<�M�<ڏ�<5��<cQ�<^��<�<�<���<��<�`�<���<��<���<�`�<��<���<�<�<^��<cQ�<5��<ڏ�<�M�<C$�<`   `   �!�<�-�<eR�<؋�<a��<�3�<p��<���<�b�<��<2��<(�<�6�<(�<2��<��<�b�<���<p��<�3�<a��<؋�<eR�<�-�<`   `   �C�<N�<�l�<��<S��<�*�<�<��<P)�<Er�<��<.��<i��<.��<��<Er�<P)�<��<�<�*�<S��<��<�l�<N�<`   `   <�<݆�<Ξ�<N��<��<�6�<,z�<���<^�<K=�<�k�<U��<�<U��<�k�<K=�<^�<���<,z�<�6�<��<N��<Ξ�<݆�<`   `   ���<X��<���<��<�+�<=X�<9��<��<���<H�<�?�<�U�<a\�<�U�<�?�<H�<���<��<9��<=X�<�+�<��<���<X��<`   `   �>�<B�<�K�<g\�<6s�<Ǝ�<���<���<Z��<��<�$�<�3�<C8�<�3�<�$�<��<Z��<���<���<Ǝ�<6s�<g\�<�K�<B�<`   `   ���<y��<���<���<���<��<���<���<" �<��<��<x �<#�<x �<��<��<" �<���<���<��<���<���<���<y��<`   `   �U�<�S�<�M�<E�<�:�<0�<�'�<Y �<J�<'�<��<�<e�<�<��<'�<J�<Y �<�'�<0�<�:�<E�<�M�<�S�<`   `   ���<���<���<��<%��<���<4u�<�X�<�A�< /�<f!�<��<��<��<f!�< /�<�A�<�X�<4u�<���<%��<��<���<���<`   `   ۣ�<���<R��<*^�<�/�<���<���<o��<*k�<NG�<�-�<�<��<�<�-�<NG�<*k�<o��<���<���<�/�<*^�<R��<���<`   `   �N�<SC�<�"�<D��<{��<�d�<��<���<���<2_�<�9�<"�<��<"�<�9�<2_�<���<���<��<�d�<{��<D��<�"�<SC�<`   `   W��<���<���<x�<�$�<��<�f�<�	�<���<�s�<�A�<�"�<��<�"�<�A�<�s�<���<�	�<�f�<��<�$�<x�<���<���<`   `   ̅�<>t�<kA�<���<Ѝ�<��<��<v7�<���<_��<aB�<��<��<��<aB�<_��<���<v7�<��<��<Ѝ�<���<kA�<>t�<`   `   9�<7��<���<FW�<���<g`�<���<zV�<���<��<�8�<�<-��<�<�8�<��<���<zV�<���<g`�<���<FW�<���<7��<`   `   ^�<uG�<��<��<��<q��<!��<�d�<?��<�u�<�$�<^��<=��<^��<�$�<�u�<?��<�d�<!��<q��<��<��<��<uG�<`   `   X��<�~�<�8�<���<�>�<��<S��<�_�<(��<R\�<��<��<t��<��<��<R\�<(��<�_�<S��<��<�>�<���<�8�<�~�<`   `   "��<���<�F�<=��<O@�<)��<���<8G�<|��<,5�<���<���<��<���<���<,5�<|��<8G�<���<)��<O@�<=��<�F�<���<`   `   ���<�|�<�0�<;��<x#�<	y�<���<��<��<��<R��<�h�<}T�<�h�<R��<��<��<��<���<	y�<x#�<;��<�0�<�|�<`   `   d_�<nE�<���<��<���<A�<��<��<�H�<M��<g�<i,�<J�<i,�<g�<M��<�H�<��<��<A�<���<��<���<nE�<`   `   H
�<���<���<'2�<��<��<�G�<��<��<i��<�'�<���<_��<���<�'�<i��<��<��<�G�<��<��<'2�<���<���<`   `   #��<^��< >�<#��<�?�<s��<&��<�R�<���<7E�<!��<���<n��<���<!��<7E�<���<�R�<&��<s��<�?�<#��< >�<^��<`   `   !"�<�
�<���<�^�<e��<@�<��<^�<W{�<i�<���< z�<�h�< z�<���<i�<W{�<^�<��<@�<e��<�^�<���<�
�<`   `   %��<���<�K�<���<Qn�<m��<GN�<	��<�=�<���<q��<�M�<[=�<�M�<q��<���<�=�<	��<GN�<m��<Qn�<���<�K�<���<`   `   ��<
�<���<�y�<%	�<\��<W�<*��<!�<p��<�^�<�/�<� �<�/�<�^�<p��<!�<*��<W�<\��<%	�<�y�<���<
�<`   `   ��<���<�`�<��<���<�<�<^��<cQ�<5��<ڏ�<�M�<C$�<��<C$�<�M�<ڏ�<5��<cQ�<^��<�<�<���<��<�`�<���<`   `   �6�<(�<2��<��<�b�<���<p��<�3�<a��<؋�<eR�<�-�<�!�<�-�<eR�<؋�<a��<�3�<p��<���<�b�<��<2��<(�<`   `   h��<.��<��<Er�<P)�<��<�<�*�<S��<��<�l�<N�<�C�<N�<�l�<��<S��<�*�<�<��<P)�<Er�<��<.��<`   `   �<U��<�k�<K=�<^�<���<,z�<�6�<��<N��<Ξ�<݆�<<�<݆�<Ξ�<N��<��<�6�<,z�<���<^�<K=�<�k�<U��<`   `   a\�<�U�<�?�<H�<���<��<9��<=X�<�+�<��<���<X��<���<X��<���<��<�+�<=X�<9��<��<���<H�<�?�<�U�<`   `   C8�<�3�<�$�<��<Z��<���<���<Ǝ�<6s�<g\�<�K�<B�<�>�<B�<�K�<g\�<6s�<Ǝ�<���<���<Z��<��<�$�<�3�<`   `   #�<x �<��<��<" �<���<���<��<���<���<���<y��<���<y��<���<���<���<��<���<���<" �<��<��<x �<`   `   e�<�<��<'�<J�<Y �<�'�<0�<�:�<E�<�M�<�S�<�U�<�S�<�M�<E�<�:�<0�<�'�<Y �<J�<'�<��<�<`   `   ��<��<f!�< /�<�A�<�X�<4u�<���<%��<��<���<���<���<���<���<��<%��<���<4u�<�X�<�A�< /�<f!�<��<`   `   ��<�<�-�<NG�<*k�<o��<���<���<�/�<*^�<R��<���<ۣ�<���<R��<*^�<�/�<���<���<o��<*k�<NG�<�-�<�<`   `   ��<"�<�9�<2_�<���<���<��<�d�<{��<D��<�"�<SC�<�N�<SC�<�"�<D��<{��<�d�<��<���<���<2_�<�9�<"�<`   `   ��<�"�<�A�<�s�<���<�	�<�f�<��<�$�<x�<���<���<W��<���<���<x�<�$�<��<�f�<�	�<���<�s�<�A�<�"�<`   `   ��<��<aB�<_��<���<v7�<��<��<Ѝ�<���<kA�<>t�<̅�<>t�<kA�<���<Ѝ�<��<��<v7�<���<_��<aB�<��<`   `   -��<�<�8�<��<���<zV�<���<g`�<���<FW�<���<7��<9�<7��<���<FW�<���<g`�<���<zV�<���<��<�8�<�<`   `   =��<^��<�$�<�u�<?��<�d�<!��<q��<��<��<��<vG�<^�<vG�<��<��<��<q��<!��<�d�<?��<�u�<�$�<^��<`   `   t��<��<��<R\�<(��<�_�<S��<��<�>�<���<�8�<�~�<X��<�~�<�8�<���<�>�<��<S��<�_�<(��<R\�<��<��<`   `   ��<���<���<,5�<|��<8G�<���<)��<P@�<=��<�F�<���<"��<���<�F�<=��<O@�<)��<���<8G�<|��<,5�<���<���<`   `   }T�<�h�<R��<��<��<��<���<	y�<x#�<;��<�0�<�|�<���<�|�<�0�<;��<x#�<	y�<���<��<��<��<R��<�h�<`   `   J�<i,�<g�<M��<�H�<��<��<A�<���<��<���<nE�<d_�<nE�<���<��<���<A�<��<��<�H�<M��<g�<i,�<`   `   _��<���<�'�<i��<��<��<�G�<��<��<'2�<���<���<H
�<���<���<'2�<��<��<�G�<��<��<i��<�'�<���<`   `   n��<���<!��<7E�<���<�R�<&��<s��<�?�<#��< >�<^��<#��<^��< >�<#��<�?�<s��<&��<�R�<���<7E�<!��<���<`   `   �h�< z�<���<i�<W{�<_�<��<@�<e��<�^�<���<�
�<!"�<�
�<���<�^�<e��<@�<��<_�<W{�<i�<���< z�<`   `   [=�<�M�<q��<���<�=�<	��<GN�<m��<Qn�<���<�K�<���<%��<���<�K�<���<Qn�<m��<GN�<	��<�=�<���<q��<�M�<`   `   � �<�/�<�^�<p��<!�<*��<W�<\��<&	�<�y�<���<
�<��<
�<���<�y�<%	�<\��<W�<*��<!�<p��<�^�<�/�<`   `   ��<L��<���<C�<�`�<<��<@�<`�<&��< ��<�8�<�]�<�i�<�]�<�8�< ��<&��<`�<@�<<��<�`�<C�<���<L��<`   `   ���<���<���<��<;T�<���<���<�2�<T|�<h��<���<�<��<�<���<h��<T|�<�2�<���<���<;T�<��<���<���<`   `   ���<��<��<�&�<�W�<��<���<��<�P�<���<Ű�<���<���<���<Ű�<���<�P�<��<���<��<�W�<�&�<��<��<`   `   t�<�<Q(�<�E�<�l�<���<[��<_�</3�<�^�<���<���<��<���<���<�^�</3�<_�<[��<���<�l�<�E�<Q(�<�<`   `   �O�<:T�<ja�<�v�<ƒ�<1��<���<S �<�$�<fE�<S^�<4n�<�t�<4n�<S^�<fE�<�$�<R �<���<1��<ƒ�<�v�<ja�<:T�<`   `   S��<��<��<I��<4��<4��<I��<��<:#�<�8�<LI�<�S�<X�<�S�<LI�<�8�<:#�<��<I��<4��<4��<I��<��<��<`   `   ��<e�<{�<��<�<L�<��<\%�<�.�<8�<@�<*E�<�F�<*E�<@�<8�<�.�<\%�<��<L�<�<��<{�<e�<`   `   1s�<@q�<Om�<-f�<�^�<�V�<�N�<"I�<~D�<�A�<�?�<?�<�=�<?�<�?�<�A�<~D�<"I�<�N�<�V�<�^�<-f�<Om�<@q�<`   `   f��< ��<���<���<߷�<I��<���<=s�<�_�<{P�<�E�<�>�<<�<�>�<�E�<{P�<�_�<=s�<���<I��<߷�<���<���< ��<`   `   �j�<ed�<S�<�7�<h�<U��<���<Π�<�~�<Xc�<O�<�B�<>�<�B�<O�<Xc�<�~�<Π�<���<U��<h�<�7�<S�<ed�<`   `   ���<���<���<��<)r�<<�<i�<m��<s��<{v�<|X�<FF�<@�<FF�<|X�<{v�<s��<m��<i�<<�<)r�<��<���<���<`   `   3_�<:U�<U6�<��<��<���<s=�<���<̹�<��<�^�<_G�<�?�<_G�<�^�<��<̹�<���<s=�<���<��<��<U6�<:U�<`   `   ���<=��<��<`�<;�<\��<Jm�<��<z��<���<�`�<�C�<�9�<�C�<�`�<���<z��<��<Jm�<\��<;�<`�<��<=��<`   `   �#�<�<���<&��<U�<��<���<�1�<&��<Z��<[�<�8�<�,�<�8�<[�<Z��<&��<�1�<���<��<U�<&��<���<�<`   `   pf�<V�<�'�<o��<���<��<���<�;�<_��<��<{L�<�&�<b�<�&�<{L�<��<_��<�;�<���<��<���<o��<�'�<V�<`   `   P��<�}�<�K�<���<N��<�$�<٬�<8�<���<�v�<�4�<�<���<�<�4�<�v�<���<8�<٬�<�$�<N��<���<�K�<�}�<`   `   ���<���<�U�<d�<��<!�<:��<�&�<s��<�Z�<��<$��<���<$��<��<�Z�<s��<�&�<:��<!�<��<d�<�U�<���<`   `   ڎ�<|�<�E�<���<���<�<���<l�<���<5�<m��<y��<F��<y��<m��<5�<���<l�<���<�<���<���<�E�<|�<`   `   �g�<�T�<W�<���<�Z�<���<P[�<V��<i�<��<k��</��<���</��<k��<��<i�<V��<P[�<���<�Z�<���<W�<�T�<`   `   �*�<��<f��<3��<�!�<A��<P&�<��<�7�<���<���<�c�<�T�<�c�<���<���<�7�<��<P&�<A��<�!�<3��<f��<��<`   `   8��<��<v��<lE�<h��<�f�<M��<Aq�<:�<Ϧ�<7a�<�5�<3'�<�5�<7a�<Ϧ�<:�<Aq�<M��<�f�<h��<lE�<v��<��<`   `   Q��<�q�<�@�<���<n��<� �<��<y8�<~��<jw�<�5�<<�<1��<<�<�5�<jw�<~��<y8�<��<� �<n��<���<�@�<�q�<`   `   #�<�<���<��<�C�<
��<mm�<��<Ԡ�<�N�<��<���<���<���<��<�N�<Ԡ�<��<mm�<
��<�C�<��<���<�<`   `   ��<��<��<L�<��<���<�5�<r��<�z�<0�<s��<���<���<���<s��<0�<�z�<r��<�5�<���<��<L�<��<��<`   `   �i�<�]�<�8�< ��<&��<`�<@�<<��<�`�<C�<���<L��<��<L��<���<C�<�`�<<��<@�<`�<&��< ��<�8�<�]�<`   `   ��<�<���<h��<T|�<�2�<���<���<;T�<��<���<���<���<���<���<��<;T�<���<���<�2�<T|�<h��<���<�<`   `   ���<���<Ű�<���<�P�<��<���<��<�W�<�&�<��<��<���<��<��<�&�<�W�<��<���<��<�P�<���<Ű�<���<`   `   ��<���<���<�^�</3�<_�<[��<���<�l�<�E�<Q(�<�<t�<�<Q(�<�E�<�l�<���<[��<_�</3�<�^�<���<���<`   `   �t�<4n�<S^�<fE�<�$�<R �<���<1��<ƒ�<�v�<ja�<:T�<�O�<:T�<ja�<�v�<ƒ�<1��<���<R �<�$�<fE�<S^�<4n�<`   `   X�<�S�<LI�<�8�<:#�<��<I��<4��<4��<I��<��<��<S��<��<��<I��<4��<4��<I��<��<:#�<�8�<KI�<�S�<`   `   �F�<*E�<@�<8�<�.�<\%�<��<L�<�<��<{�<e�<��<e�<{�<��<�<L�<��<\%�<�.�<8�<@�<*E�<`   `   �=�<?�<�?�<�A�<~D�<"I�<�N�<�V�<�^�<-f�<Om�<@q�<1s�<@q�<Om�<-f�<�^�<�V�<�N�<"I�<~D�<�A�<�?�<?�<`   `   <�<�>�<�E�<{P�<�_�<=s�<���<I��<߷�<���<���< ��<f��< ��<���<���<߷�<I��<���<=s�<�_�<{P�<�E�<�>�<`   `   >�<�B�<O�<Xc�<�~�<Π�<���<U��<h�<�7�<S�<ed�<�j�<ed�<S�<�7�<h�<U��<���<Π�<�~�<Xc�<O�<�B�<`   `   @�<FF�<|X�<{v�<s��<m��<i�<<�<)r�<��<���<���<���<���<���<��<)r�<<�<i�<m��<s��<{v�<|X�<FF�<`   `   �?�<_G�<�^�<��<̹�<���<s=�<���<��<��<U6�<:U�<3_�<:U�<U6�<��<��<���<s=�<���<̹�<��<�^�<_G�<`   `   �9�<�C�<�`�<���<z��<��<Jm�<\��<;�<`�<��<=��<���<=��<��<`�<;�<\��<Jm�<��<z��<���<�`�<�C�<`   `   �,�<�8�<[�<Z��<&��<�1�<���<��<U�<&��<���<�<�#�<�<���<&��<U�<��<���<�1�<&��<Z��<[�<�8�<`   `   b�<�&�<{L�<��<`��<�;�<���<��<���<o��<�'�<V�<pf�<V�<�'�<o��<���<��<���<�;�<_��<��<{L�<�&�<`   `   ���<�<�4�<�v�<���<8�<٬�<�$�<N��<���<�K�<�}�<P��<�}�<�K�<���<N��<�$�<٬�<8�<���<�v�<�4�<�<`   `   ���<$��<��<�Z�<s��<�&�<:��<!�<��<d�<�U�<���<���<���<�U�<d�<��<!�<:��<�&�<s��<�Z�<��<$��<`   `   F��<y��<m��<5�<���<l�<���<�<���<���<�E�<|�<ڎ�<|�<�E�<���<���<�<���<l�<���<5�<m��<y��<`   `   ���</��<k��<��<i�<V��<P[�<���<�Z�<���<W�<�T�<�g�<�T�<W�<���<�Z�<���<P[�<V��<i�<��<k��</��<`   `   �T�<�c�<���<���<�7�<��<P&�<A��<�!�<3��<g��<��<�*�<��<f��<3��<�!�<A��<P&�<��<�7�<���<���<�c�<`   `   3'�<�5�<7a�<Ϧ�<:�<Aq�<M��<�f�<h��<lE�<v��<��<8��<��<v��<lE�<h��<�f�<M��<Aq�<:�<Ϧ�<7a�<�5�<`   `   1��<<�<�5�<jw�<~��<y8�<��<� �<n��<���<�@�<�q�<Q��<�q�<�@�<���<n��<� �<��<y8�<~��<jw�<�5�<<�<`   `   ���<���<��<�N�<Ԡ�<��<mm�<
��<�C�<��<���<�<#�<�<���<��<�C�<
��<mm�<��<Ԡ�<�N�<��<���<`   `   ���<���<s��<0�<�z�<r��<�5�<���<��<L�<��<��<��<��<��<L�<��<���<�5�<r��<�z�<0�<s��<���<`   `   \?�<H�<"`�<���<��<���<T6�<�x�<��<M��<��<�4�<.>�<�4�<��<M��<��<�x�<T6�<���<��<���<"`�<H�<`   `   %F�<�M�<�a�<���<���</��<��<�V�<���<]��<���<+��<�<+��<���<]��<���<�V�<��</��<���<���<�a�<�M�<`   `   #Z�<v`�<.q�<���<���<���<	�<�>�<�l�<���<��<���<o��<���<��<���<�l�<�>�<	�<���<���<���<.q�<v`�<`   `   �{�<2��<��<J��<���<���<�<�0�<4V�<�v�<���<��<��<��<���<�v�<4V�<�0�<�<���<���<J��<��<2��<`   `   ���<��<Ϲ�<(��<��<K��<��<�/�<�J�<�b�<Nu�<���<���<���<Nu�<�b�<�J�<�/�<��<K��<��<(��<Ϲ�<��<`   `   ���<��<���<���<3�<��<�&�<�8�<-J�<Y�<�d�<yl�<4o�<yl�<�d�<Y�<-J�<�8�<�&�<��<3�<���<���<��<`   `   `4�<4�<�5�<�7�<#;�<�?�<�D�<|K�<PR�<(X�<-]�<�`�<�a�<�`�<-]�<(X�<PR�<|K�<�D�<�?�<#;�<�7�<�5�<4�<`   `   ׇ�<��<Ղ�<o}�<qw�<hq�<#k�<�e�<�a�<�^�<�\�<)\�<�[�<)\�<�\�<�^�<�a�<�e�<#k�<hq�<qw�<o}�<Ղ�<��<`   `   ���<n��<���<���<���<a��<n��<���<5v�<Wj�<a�<�[�<[Z�<�[�<a�<Wj�<5v�<���<n��<a��<���<���<���<n��<`   `   l>�<�9�<\-�<	�<���<���<���<���<���<�x�<>h�<f^�<�[�<f^�<>h�<�x�<���<���<���<���<���<	�<\-�<�9�<`   `   ���<��<��<�f�<D�<3�<r��<���<(��<��<�o�<�a�<]�<�a�<�o�<��<(��<���<r��<3�<D�<�f�<��<��<`   `   ���<���<��<���<P��<�Q�<��<���<���<���<Nu�<�b�<�\�<�b�<Nu�<���<���<���<��<�Q�<P��<���<��<���<`   `   +?�<�6�<X�<���<��<`��<�@�<C�<���<N��<�v�<�`�<UY�<�`�<�v�<N��<���<C�<�@�<`��<��<���<X�<�6�<`   `   8��<�u�<�W�<�'�<1��<��<�[�<�<��<T��<9s�<�Y�<�Q�<�Y�<9s�<T��<��<�<�[�<��<1��<�'�<�W�<�u�<`   `   ��<���<7��<)N�<
�<ɼ�<Bk�<#�<���<���<�h�<=L�<C�<=L�<�h�<���<���<#�<Bk�<ɼ�<
�<)N�<7��<���<`   `   ���<v��<:��<9d�<�<,��<o�<��<'��<K��<�W�<^8�<.�<^8�<�W�<K��<'��<��<o�<,��<�<9d�<:��<v��<`   `   ��<~��<s��<Th�<��<2��<cf�<O�<ع�<lt�<�?�<\�<��<\�<�?�<lt�<ع�<O�<cf�<2��<��<Th�<s��<~��<`   `   n��<Q��<��<[�<:�<���<FR�<N��<��<HX�<u"�<+�<.��<+�<u"�<HX�<��<N��<FR�<���<:�<[�<��<Q��<`   `   c��<ѣ�<6|�<�=�<���<���<�3�<���<��<g7�<� �<���<w��<���<� �<g7�<��<���<�3�<���<���<�=�<6|�<ѣ�<`   `   ��<�w�<�P�<��<��<�j�<9�<~��<sZ�<#�<���<-��<���<-��<���<#�<sZ�<~��<9�<�j�<��<��<�P�<�w�<`   `   LL�<�?�<s�<(��<��<|;�<���<܅�<:3�<���<��<!��<@��<!��<��<���<:3�<܅�<���<|;�<��<(��<s�<�?�<`   `   ?�<\��<���<N��<,[�<a�<��<�[�<8�<���<���<�y�<|n�<�y�<���<���<8�<�[�<��<a�<,[�<N��<���<\��<`   `   E��<ɺ�<<��<�d�<�!�<���<��<�2�<���<ɫ�<
}�<A`�<HV�<A`�<
}�<ɫ�<���<�2�<��<���<�!�<�d�<<��<ɺ�<`   `   ���<v�<�W�<�'�<���<��<CY�<��<���<p��<Ti�<�N�<�E�<�N�<Ti�<p��<���<��<CY�<��<���<�'�<�W�<v�<`   `   .>�<�4�<��<M��<��<�x�<T6�<���<��<���<"`�<H�<\?�<H�<"`�<���<��<���<T6�<�x�<��<M��<��<�4�<`   `   �<+��<���<]��<���<�V�<��</��<���<���<�a�<�M�<%F�<�M�<�a�<���<���</��<��<�V�<���<]��<���<+��<`   `   o��<���<��<���<�l�<�>�<	�<���<���<���<.q�<v`�<#Z�<v`�<.q�<���<���<���<	�<�>�<�l�<���<��<���<`   `   ��<��<���<�v�<4V�<�0�<�<���<���<J��<��<2��<�{�<2��<��<J��<���<���<�<�0�<4V�<�v�<���<��<`   `   ���<���<Nu�<�b�<�J�<�/�<��<K��<��<(��<ι�<��<���<��<ι�<(��<��<K��<��<�/�<�J�<�b�<Nu�<���<`   `   4o�<yl�<�d�<Y�<-J�<�8�<�&�<��<3�<���<���<��<���<��<���<���<3�<��<�&�<�8�<-J�<Y�<�d�<yl�<`   `   �a�<�`�<-]�<(X�<PR�<|K�<�D�<�?�<#;�<�7�<�5�<4�<`4�<4�<�5�<�7�<#;�<�?�<�D�<|K�<PR�<(X�<-]�<�`�<`   `   �[�<)\�<�\�<�^�<�a�<�e�<#k�<hq�<qw�<o}�<Ղ�<��<ׇ�<��<Ղ�<o}�<qw�<hq�<#k�<�e�<�a�<�^�<�\�<)\�<`   `   [Z�<�[�<a�<Wj�<5v�<���<n��<a��<���<���<���<n��<���<n��<���<���<���<a��<n��<���<5v�<Wj�<a�<�[�<`   `   �[�<f^�<>h�<�x�<���<���<���<���<���<	�<\-�<�9�<l>�<�9�<\-�<	�<���<���<���<���<���<�x�<>h�<f^�<`   `   ]�<�a�<�o�<��<(��<���<r��<3�<D�<�f�<��<��<���<��<��<�f�<D�<3�<r��<���<(��<��<�o�<�a�<`   `   �\�<�b�<Nu�<���<���<���<��<�Q�<P��<���<��<���<���<���<��<���<P��<�Q�<��<���<���<���<Nu�<�b�<`   `   UY�<�`�<�v�<N��<���<C�<�@�<`��<��<���<X�<�6�<+?�<�6�<X�<���<��<`��<�@�<C�<���<N��<�v�<�`�<`   `   �Q�<�Y�<9s�<T��<��<�<�[�<��<1��<�'�<�W�<�u�<8��<�u�<�W�<�'�<1��<��<�[�<�<��<T��<9s�<�Y�<`   `   C�<=L�<�h�<���<���<#�<Bk�<ɼ�<
�<)N�<7��<���<��<���<7��<)N�<
�<ɼ�<Bk�<#�<���<���<�h�<=L�<`   `   .�<^8�<�W�<K��<'��<��<o�<,��<�<9d�<:��<v��<���<v��<:��<9d�<�<,��<o�<��<'��<K��<�W�<^8�<`   `   ��<\�<�?�<lt�<ع�<O�<cf�<2��<��<Th�<s��<~��<��<~��<s��<Th�<��<2��<cf�<O�<ع�<lt�<�?�<\�<`   `   .��<+�<u"�<HX�<��<N��<FR�<���<:�<[�<��<Q��<n��<Q��<��<[�<:�<���<FR�<N��<��<HX�<u"�<+�<`   `   w��<���<� �<g7�<��<���<�3�<���<���<�=�<6|�<ѣ�<c��<ѣ�<6|�<�=�<���<���<�3�<���<��<g7�<� �<���<`   `   ���<-��<���<#�<sZ�<~��<9�<�j�<��<��<�P�<�w�<��<�w�<�P�<��<��<�j�<9�<~��<sZ�<#�<���<-��<`   `   @��<!��<��<���<:3�<܅�<���<|;�<��<(��<s�<�?�<LL�<�?�<s�<(��<��<|;�<���<܅�<:3�<���<��<!��<`   `   |n�<�y�<���<���<9�<�[�<��<a�<,[�<N��<���<\��<?�<\��<���<N��<,[�<a�<��<�[�<8�<���<���<�y�<`   `   HV�<A`�<
}�<ɫ�<���<�2�<��<���<�!�<�d�<<��<ɺ�<F��<ɺ�<<��<�d�<�!�<���<��<�2�<���<ɫ�<
}�<A`�<`   `   �E�<�N�<Ti�<p��<���<��<CY�<��<���<�'�<�W�<v�<���<v�<�W�<�'�<���<��<CY�<��<���<p��<Ti�<�N�<`   `   ���<���<b��<��<)��<�'�<�X�<��<���<w��<�<��<)�<��<�<w��<���<��<�X�<�'�<)��<��<b��<���<`   `   ���</��<޸�<���<)��<��<�D�<�o�<��<k��<���<���<L��<���<���<k��<��<�o�<�D�<��<)��<���<޸�</��<`   `   ��<|��<f��<���<K��<`�<�9�<�]�<6��<۝�<8��<���<��<���<8��<۝�<6��<�]�<�9�<`�<K��<���<f��<|��<`   `   M��<��<S��<��<� �<��<7�<wT�<�o�<���<Ù�<p��<,��<p��<Ù�<���<�o�<wT�<7�<��<� �<��<S��<��<`   `    ��<���<���<��<��<�(�<=�<�R�<�f�<Rw�<߅�<���<ΐ�<���<߅�<Rw�<�f�<�R�<=�<�(�<��<��<���<���<`   `   r�<� �<�$�<Y,�<X5�<@�<�L�<uY�<�e�<Qp�<�y�<�<I��<�<�y�<Qp�<�e�<uY�<�L�<@�<X5�<Y,�<�$�<� �<`   `   �U�<jV�<�W�<�Y�<m[�<�^�<kc�<9g�<�k�<�o�<Bs�<|u�<v�<|u�<Bs�<�o�<�k�<9g�<kc�<�^�<m[�<�Y�<�W�<jV�<`   `   ��<���<��<v��<���<���<�<z�<�v�<�t�<jr�<wq�<Fq�<wq�<jr�<�t�<�v�<z�<�<���<���<v��<��<���<`   `   ,��<<��<��<���<*��<Ӭ�<��<��<ۆ�<v}�<v�<�q�< p�<�q�<v�<v}�<ۆ�<��<��<Ӭ�<*��<���<��<<��<`   `   
�<��<S�<g �<w��<��<���<��<S��<���<2{�<�s�<�p�<�s�<2{�<���<S��<��<���<��<w��<g �<S�<��<`   `   i`�<�[�<�N�<;�<� �<��<p��<S��<���<��<��<&v�<`r�<&v�<��<��<���<S��<p��<��<� �<;�<�N�<�[�<`   `   f��<a��<"��<q�<�O�<R*�<��<���<���<���<��<�w�<�r�<�w�<��<���<���<���<��<R*�<�O�<q�<"��<a��<`   `   M��<M��<Ⱦ�<���<Fy�<M�<��<���<t��<ա�<F��<)v�<}p�<)v�<F��<ա�<t��<���<��<M�<Fy�<���<Ⱦ�<M��<`   `   U�<� �<���<���<��<h�<x1�<-��<��<M��<��<�p�<�j�<�p�<��<M��<��<-��<x1�<h�<��<���<���<� �<`   `   �*�<�"�<B
�<��<f��<+y�<!=�<w�<���<��<�|�<�g�<�`�<�g�<�|�<��<���<w�<!=�<+y�<f��<��<B
�<�"�<`   `   �@�<�7�<��<���<\��<��<�@�<�<���<���<�p�<�Y�<�Q�<�Y�<�p�<���<���<�<�@�<��<\��<���<��<�7�<`   `   �G�<Q>�<S"�<���<S��<1~�<n:�<��<���<
��<_�<�F�<�=�<�F�<_�<
��<���<��<n:�<1~�<S��<���<S"�<Q>�<`   `   i@�<�6�<4�<O��<���<�p�<�*�<���<��<�q�<I�<�/�<'�<�/�<I�<�q�<��<���<�*�<�p�<���<O��<4�<�6�<`   `   �+�<�!�<g�<H��<ԝ�<�Z�<��<s��<��<GY�<�0�<��<��<��<�0�<GY�<��<s��<��<�Z�<ԝ�<H��<g�<�!�<`   `   ��<	�<���<��<��<5=�<E��<s��</s�<>�<��<N��<���<N��<��<>�</s�<s��<E��<5=�<��<��<���<	�<`   `   ���<a��<n��<��<VZ�<�<G��< ��<�U�<"�<k��<���<���<���<k��<"�<�U�< ��<G��<�<VZ�<��<n��<a��<`   `   8��<1��<��<�f�<K1�<��<���<'s�<89�<��<���<p��<=��<p��<���<��<89�<'s�<���<��<K1�<�f�<��<1��<`   `   1��<�w�<�_�<_9�<��<���<c��<qU�<$�<���<��<U��<Я�<U��<��<���<$�<qU�<c��<���<��<_9�<�_�<�w�<`   `   ZM�<6E�</�<��<���<���<_r�<�;�<j	�<���<N��<@��<c��<@��<N��<���<j	�<�;�<_r�<���<���<��</�<6E�<`   `   )�<��<�<w��<���<��<�X�<�'�<)��<��<b��<���<���<���<b��<��<)��<�'�<�X�<��<���<w��<�<��<`   `   L��<���<���<k��<��<�o�<�D�<��<)��<���<޸�</��<���</��<޸�<���<)��<��<�D�<�o�<��<k��<���<���<`   `   ��<���<8��<۝�<6��<�]�<�9�<`�<K��<���<f��<|��<��<|��<f��<���<K��<`�<�9�<�]�<6��<۝�<8��<���<`   `   ,��<p��<Ù�<���<�o�<wT�<7�<��<� �<��<S��<��<M��<��<S��<��<� �<��<7�<wT�<�o�<���<Ù�<p��<`   `   ΐ�<���<߅�<Rw�<�f�<�R�<=�<�(�<��<��<���<���< ��<���<���<��<��<�(�<=�<�R�<�f�<Rw�<߅�<���<`   `   I��<�<�y�<Qp�<�e�<uY�<�L�<@�<X5�<Y,�<�$�<� �<r�<� �<�$�<Y,�<X5�<@�<�L�<uY�<�e�<Qp�<�y�<�<`   `   v�<|u�<Bs�<�o�<�k�<9g�<kc�<�^�<m[�<�Y�<�W�<jV�<�U�<jV�<�W�<�Y�<m[�<�^�<kc�<9g�<�k�<�o�<Bs�<|u�<`   `   Fq�<wq�<jr�<�t�<�v�<z�<�<���<���<v��<��<���<��<���<��<v��<���<���<�<z�<�v�<�t�<jr�<wq�<`   `    p�<�q�<v�<v}�<ۆ�<��<��<Ӭ�<*��<���<��<<��<,��<<��<��<���<*��<Ӭ�<��<��<ۆ�<v}�<v�<�q�<`   `   �p�<�s�<2{�<���<S��<��<���<��<w��<g �<S�<��<
�<��<S�<g �<w��<��<���<��<S��<���<2{�<�s�<`   `   `r�<&v�<��<��<���<S��<p��<��<� �<;�<�N�<�[�<i`�<�[�<�N�<;�<� �<��<p��<S��<���<��<��<&v�<`   `   �r�<�w�<��<���<���<���<��<R*�<�O�<q�<"��<a��<f��<a��<"��<q�<�O�<R*�<��<���<���<���<��<�w�<`   `   }p�<)v�<F��<ա�<t��<���<��<M�<Fy�<���<Ⱦ�<M��<M��<M��<Ⱦ�<���<Fy�<M�<��<���<t��<ա�<F��<)v�<`   `   �j�<�p�<��<M��<��<-��<x1�<h�<��<���<���<� �<U�<� �<���<���<��<h�<x1�<-��<��<M��<��<�p�<`   `   �`�<�g�<�|�<��<���<w�<!=�<+y�<f��<��<B
�<�"�<�*�<�"�<B
�<��<f��<+y�<!=�<w�<���<��<�|�<�g�<`   `   �Q�<�Y�<�p�<���<���<�<�@�<��<\��<���<��<�7�<�@�<�7�<��<���<\��<��<�@�<�<���<���<�p�<�Y�<`   `   �=�<�F�<_�<
��<���<��<n:�<1~�<S��<���<S"�<Q>�<�G�<Q>�<S"�<���<S��<1~�<n:�<��<���<
��<_�<�F�<`   `   '�<�/�<I�<�q�<��<���<�*�<�p�<���<O��<4�<�6�<i@�<�6�<4�<O��<���<�p�<�*�<���<��<�q�<I�<�/�<`   `   ��<��<�0�<GY�<��<s��<��<�Z�<ԝ�<H��<g�<�!�<�+�<�!�<g�<H��<ԝ�<�Z�<��<s��<��<GY�<�0�<��<`   `   ���<N��<��<>�</s�<s��<E��<5=�<��<��<���<	�<��<	�<���<��<��<5=�<E��<s��</s�<>�<��<N��<`   `   ���<���<k��<"�<�U�< ��<G��<�<VZ�<��<n��<a��<���<a��<n��<��<VZ�<�<G��< ��<�U�<"�<k��<���<`   `   =��<p��<���<��<89�<'s�<���<��<K1�<�f�<��<1��<8��<1��<��<�f�<K1�<��<���<'s�<89�<��<���<p��<`   `   Я�<U��<��<���<$�<qU�<c��<���<��<_9�<�_�<�w�<1��<�w�<�_�<_9�<��<���<c��<qU�<$�<���<��<U��<`   `   c��<@��<N��<���<j	�<�;�<_r�<���<���<��</�<6E�<ZM�<6E�</�<��<���<���<_r�<�;�<j	�<���<N��<@��<`   `   U��<&��<���<��<�)�<yK�<�o�<ɕ�<v��<��<���<���<f�<���<���<��<v��<ɕ�<�o�<yK�<�)�<��<���<&��<`   `   f��<���<���<�<�$�<B�<�a�<U��<���<��<Q��<��<���<��<Q��<��<���<U��<�a�<B�<�$�<�<���<���<`   `   ���<���<
�<��</&�< ?�<zY�<_t�<���<F��<"��<��<���<��<"��<F��<���<_t�<zY�< ?�</&�<��<
�<���<`   `   �<�
�<S�<��</�<�B�<�W�<Rm�<>��<<��<m��<��<"��<��<m��<<��<>��<Rm�<�W�<�B�</�<��<S�<�
�<`   `   �"�<�$�<l*�<a3�<c?�<M�<f\�<�k�<�z�<ˇ�<[��<���<
��<���<[��<ˇ�<�z�<�k�<f\�<M�<c?�<a3�<l*�<�$�<`   `   wE�<
G�<�I�<�N�<�U�<W^�<�g�<Jp�<ry�<ہ�<���<���<���<���<���<ہ�<ry�<Jp�<�g�<W^�<�U�<�N�<�I�<
G�<`   `   �n�<�o�<�o�<�p�<�r�<�t�<�w�<�z�<
~�<.��<O��<���<Ӆ�<���<O��<.��<
~�<�z�<�w�<�t�<�r�<�p�<�o�<�o�<`   `   ��<��<���<���<˔�<���<���<���<͆�<2��<ނ�<ā�<���<ā�<ނ�<2��<͆�<���<���<���<˔�<���<���<��<`   `   ���<���<���<A��<���<y��<��<?��<(��<��<=��<́�<6��<́�<=��<��<(��<?��<��<y��<���<A��<���<���<`   `   ��<u��<m��<s��<��<H��<���<׭�<��<p��<���<���<@��<���<���<p��<��<׭�<���<H��<��<s��<m��<u��<`   `   �3�<�0�<)'�<�<��<��<���<���<Z��<��<���<L��<���<L��<���<��<Z��<���<���<��<��<�<)'�<�0�<`   `   �b�<�^�<�R�<@�<(�<��<8��<n��<��<��<���<?��<B��<?��<���<��<��<n��<8��<��<(�<@�<�R�<�^�<`   `   ���<ȇ�<�y�<Kc�<�F�<^%�<��<���<���<L��<<��<Ӆ�<���<Ӆ�<<��<L��<���<���<��<^%�<�F�<Kc�<�y�<ȇ�<`   `   ���<s��<9��<��<_�<9�<��<���<i��<٧�<���<q��<}�<q��<���<٧�<i��<���<��<9�<_�<��<9��<s��<`   `   ���<T��<u��<9��<+p�<fF�<��<��<"��</��<x��<a{�<�u�<a{�<x��</��<"��<��<��<fF�<+p�<9��<u��<T��<`   `   ���<���<[��<��<�x�<�K�<k�<6��<m��<ݝ�<���<�p�<�j�<�p�<���<ݝ�<m��<6��<k�<�K�<�x�<��<[��<���<`   `   ���<���<���<k��<$y�<�I�<��<I��<Q��<Ē�<$u�<,c�<�\�<,c�<$u�<Ē�<Q��<I��<��<�I�<$y�<k��<���<���<`   `   ���<7��<���<o��<q�<L@�<��<��<X��<{��<�d�<GR�<�K�<GR�<�d�<{��<X��<��<��<L@�<q�<o��<���<7��<`   `   ��<���<Ĭ�<���<�`�<�/�<���<d��<И�<xp�<>R�<r?�<�8�<r?�<>R�<xp�<И�<d��<���<�/�<�`�<���<Ĭ�<���<`   `   u��<u��<��<u�<�J�<��<P��<���<���<i\�<S>�<]+�<�$�<]+�<S>�<i\�<���<���<P��<��<�J�<u�<��<u��<`   `   7��<h��<mx�<�X�<�/�<. �<���<���</o�<�G�<Y*�<��<��<��<Y*�<�G�</o�<���<���<. �<�/�<�X�<mx�<h��<`   `   �p�<9j�<�V�<�8�<v�<2��<R��<���<�X�<�3�<��<w�<� �<w�<��<�3�<�X�<���<R��<2��<v�<�8�<�V�<9j�<`   `   CK�<XE�<f3�<��<~��<���<"��<�n�<QE�<�"�<e�<���<���<���<e�<�"�<QE�<�n�<"��<���<~��<��<f3�<XE�<`   `   j%�<5 �<��<7��<	��<��<\��< [�<R5�<��<O��<���<���<���<O��<��<R5�< [�<\��<��<	��<7��<��<5 �<`   `   f�<���<���<��<v��<ɕ�<�o�<yK�<�)�<��<���<&��<U��<&��<���<��<�)�<yK�<�o�<ɕ�<v��<��<���<���<`   `   ���<��<Q��<��<���<U��<�a�<B�<�$�<�<���<���<f��<���<���<�<�$�<B�<�a�<U��<���<��<Q��<��<`   `   ���<��<"��<F��<���<_t�<zY�< ?�</&�<��<
�<���<���<���<
�<��</&�< ?�<zY�<_t�<���<F��<"��<��<`   `   "��<��<m��<<��<>��<Rm�<�W�<�B�</�<��<S�<�
�<�<�
�<S�<��</�<�B�<�W�<Rm�<>��<<��<m��<��<`   `   
��<���<[��<ˇ�<�z�<�k�<f\�<M�<c?�<a3�<l*�<�$�<�"�<�$�<l*�<a3�<c?�<M�<f\�<�k�<�z�<ˇ�<[��<���<`   `   ���<���<���<ہ�<ry�<Jp�<�g�<W^�<�U�<�N�<�I�<
G�<wE�<
G�<�I�<�N�<�U�<W^�<�g�<Jp�<ry�<ہ�<���<���<`   `   Ӆ�<���<O��<.��<
~�<�z�<�w�<�t�<�r�<�p�<�o�<�o�<�n�<�o�<�o�<�p�<�r�<�t�<�w�<�z�<
~�<.��<O��<���<`   `   ���<ā�<ނ�<2��<͆�<���<���<���<˔�<���<���<��<��<��<���<���<˔�<���<���<���<͆�<2��<ނ�<ā�<`   `   6��<́�<=��<��<(��<?��<��<y��<���<A��<���<���<���<���<���<A��<���<y��<��<?��<(��<��<=��<́�<`   `   @��<���<���<p��<��<׭�<���<H��<��<s��<m��<u��<��<u��<m��<s��<��<H��<���<׭�<��<p��<���<���<`   `   ���<L��<���<��<Z��<���<���<��<��<�<)'�<�0�<�3�<�0�<)'�<�<��<��<���<���<Z��<��<���<L��<`   `   B��<?��<���<��<��<n��<8��<��<(�<@�<�R�<�^�<�b�<�^�<�R�<@�<(�<��<8��<n��<��<��<���<?��<`   `   ���<Ӆ�<<��<M��<���<���<��<^%�<�F�<Kc�<�y�<ɇ�<���<ȇ�<�y�<Kc�<�F�<^%�<��<���<���<L��<<��<Ӆ�<`   `   }�<q��<���<٧�<i��<���<��<9�<_�<��<9��<s��<���<s��<9��<��<_�<9�<��<���<i��<٧�<���<q��<`   `   �u�<a{�<x��</��<"��<��<��<fF�<+p�<9��<u��<T��<���<T��<u��<9��<+p�<fF�<��<��<"��</��<x��<a{�<`   `   �j�<�p�<���<ݝ�<m��<6��<k�<�K�<�x�<��<[��<���<���<���<[��<��<�x�<�K�<k�<6��<m��<ݝ�<���<�p�<`   `   �\�<,c�<$u�<Ē�<Q��<I��<��<�I�<$y�<k��<���<���<���<���<���<k��<$y�<�I�<��<I��<Q��<Ē�<$u�<,c�<`   `   �K�<GR�<�d�<{��<X��<��<��<L@�<q�<o��<���<7��<���<7��<���<o��<q�<L@�<��<��<X��<{��<�d�<GR�<`   `   �8�<r?�<>R�<xp�<И�<d��<���<�/�<�`�<���<Ĭ�<���<��<���<Ĭ�<���<�`�<�/�<���<d��<И�<xp�<>R�<r?�<`   `   �$�<]+�<S>�<i\�<���<���<P��<��<�J�<u�<��<u��<u��<u��<��<u�<�J�<��<P��<���<���<i\�<S>�<]+�<`   `   ��<��<Y*�<�G�</o�<���<���<. �<�/�<�X�<mx�<h��<7��<h��<mx�<�X�<�/�<. �<���<���</o�<�G�<Y*�<��<`   `   � �<w�<��<�3�<�X�<���<R��<2��<v�<�8�<�V�<9j�<�p�<9j�<�V�<�8�<v�<2��<R��<���<�X�<�3�<��<w�<`   `   ���<���<e�<�"�<QE�<�n�<"��<���<~��<��<f3�<XE�<CK�<XE�<f3�<��<~��<���<"��<�n�<QE�<�"�<e�<���<`   `   ���<���<O��<��<R5�< [�<\��<��<	��<7��<��<5 �<j%�<5 �<��<7��<	��<��<\��< [�<R5�<��<O��<���<`   `   a�<��<'�<7�<CM�<Af�<���<���<^��<>��<C��<J��<���<J��<C��<>��<^��<���<���<Af�<CM�<7�<'�<��<`   `   %�<-�<W(�<y6�<AI�<�^�<�v�<���<��<���<���<Z��<9��<Z��<���<���<��<���<�v�<�^�<AI�<y6�<W(�<-�<`   `   �$�<)'�<�.�<s:�<OJ�<G\�<Hp�<���<Q��<���<
��<a��<���<a��<
��<���<Q��<���<Hp�<G\�<OJ�<s:�<�.�<)'�<`   `   �3�<.5�<2;�<gD�<Q�<&_�<�n�<�~�<R��<Κ�<���<_��<I��<_��<���<Κ�<R��<�~�<�n�<&_�<Q�<gD�<2;�<.5�<`   `   �G�<I�<�M�<�S�<�\�<�f�<�r�<�}�<���<~��<���<z��<��<z��<���<~��<���<�}�<�r�<�f�<�\�<�S�<�M�<I�<`   `   �a�<Eb�<�d�<�h�<�m�<�s�<z�<���<?��<���<$��<���<��<���<$��<���<?��<���<z�<�s�<�m�<�h�<�d�<Eb�<`   `   `��<f��<��<S��<���<;��<Y��<��<8��<���<ێ�<���<��<���<ێ�<���<8��<��<Y��<;��<���<S��<��<f��<`   `   ���<��<���<ʞ�<��<a��<I��<���<���<���<���<j��<i��<j��<���<���<���<���<I��<a��<��<ʞ�<���<��<`   `   T��<G��<��<���<���<��<���<���<
��<4��<ُ�<+��<���<+��<ُ�<4��<
��<���<���<��<���<���<��<G��<`   `   h��<���<k��<���<���<���<B��<Ѯ�<ܣ�<i��<ْ�<x��<1��<x��<ْ�<i��<ܣ�<Ѯ�<B��<���<���<���<k��<���<`   `   =�<��<��<���<���<'��<-��<]��<���<���<h��<��< ��<��<h��<���<���<]��<-��<'��<���<���<��<��<`   `   �4�<2�<U)�<��<�	�<��<s��<���<���<��<���<'��<���<'��<���<��<���<���<s��<��<�	�<��<U)�<2�<`   `   )S�<�O�<�E�<M5�<p �<��<���<m��<'��<���<��<А�<]��<А�<��<���<'��<m��<���<��<p �<M5�<�E�<�O�<`   `   �l�<rh�<�\�<*J�<;2�<K�<���<���<��<H��<��<���<u��<���<��<H��<��<���<���<K�<;2�<*J�<�\�<rh�<`   `   ��<{�<�m�<CY�<�>�<: �<���<��<���<]��<.��<���<b��<���<.��<]��<���<��<���<: �<�>�<CY�<�m�<{�<`   `   Ҋ�<ޅ�<x�<�a�<CE�<P$�<� �<r��<���<_��<h��<v��<J}�<v��<h��<_��<���<r��<� �<P$�<CE�<�a�<x�<ޅ�<`   `   ���<p��<�z�<0c�<\E�<f"�</��<@��<��<���<2��<Zw�<�r�<Zw�<2��<���<��<@��</��<f"�<\E�<0c�<�z�<p��<`   `   ���<���<ov�<�]�<�?�<o�<@��<���<���<���<4y�<�j�<Ff�<�j�<4y�<���<���<���<@��<o�<�?�<�]�<ov�<���<`   `   ��<�z�<	k�<mR�<�3�<g�<���<���<���<��<�j�<�\�<JX�<�\�<�j�<��<���<���<���<g�<�3�<mR�<	k�<�z�<`   `   �n�<Vi�<1Z�<.B�<	#�<v��<��<���<Y��<�r�<1\�<!N�<nI�<!N�<1\�<�r�<Y��<���<��<v��<	#�<.B�<1Z�<Vi�<`   `   �X�<mS�<E�<�-�<$�<o��<���<���<��<:c�<jM�<o?�<�:�<o?�<jM�<:c�<��<���<���<o��<$�<�-�<E�<mS�<`   `   <?�<b:�<J,�<��<���<`��<y��<���<�o�<fT�<O?�<�1�<�-�<�1�<O?�<fT�<�o�<���<y��<`��<���<��<J,�<b:�<`   `   �#�<U�<��<���<���<q��<��<��<ua�<�G�<�3�<%'�<#�<%'�<�3�<�G�<ua�<��<��<q��<���<���<��<U�<`   `   ��<��<i��<p��<]��<M��<��<dq�<{U�<�=�<N+�<��<��<��<N+�<�=�<{U�<dq�<��<M��<]��<p��<i��<��<`   `   ���<J��<C��<>��<^��<���<���<Af�<CM�<7�<'�<��<a�<��<'�<7�<CM�<Af�<���<���<^��<>��<C��<J��<`   `   9��<Z��<���<���<��<���<�v�<�^�<AI�<y6�<W(�<-�<%�<-�<W(�<y6�<AI�<�^�<�v�<���<��<���<���<Z��<`   `   ���<a��<
��<���<Q��<���<Hp�<G\�<OJ�<s:�<�.�<)'�<�$�<)'�<�.�<s:�<OJ�<G\�<Hp�<���<Q��<���<
��<a��<`   `   I��<_��<���<Κ�<R��<�~�<�n�<&_�<Q�<gD�<2;�<.5�<�3�<.5�<2;�<gD�<Q�<&_�<�n�<�~�<R��<Κ�<���<_��<`   `   ��<z��<���<~��<���<�}�<�r�<�f�<�\�<�S�<�M�<I�<�G�<I�<�M�<�S�<�\�<�f�<�r�<�}�<���<~��<���<z��<`   `   ��<���<$��<���<?��<���<z�<�s�<�m�<�h�<�d�<Eb�<�a�<Eb�<�d�<�h�<�m�<�s�<z�<���<?��<���<$��<���<`   `   ��<���<ێ�<���<8��<��<Y��<;��<���<S��<��<f��<`��<f��<��<S��<���<;��<Y��<��<8��<���<ێ�<���<`   `   i��<j��<���<���<���<���<I��<a��<��<ʞ�<���<��<���<��<���<ʞ�<��<a��<I��<���<���<���<���<j��<`   `   ���<+��<ُ�<4��<
��<���<���<��<���<���<��<F��<T��<F��<��<���<���<��<���<���<
��<4��<ُ�<+��<`   `   1��<x��<ْ�<i��<ܣ�<Ѯ�<B��<���<���<���<k��<���<h��<���<k��<���<���<���<B��<Ѯ�<ܣ�<i��<ْ�<x��<`   `    ��<��<h��<���<���<]��<-��<'��<���<���<��<��<=�<��<��<���<���<'��<-��<]��<���<���<h��<��<`   `   ���<'��<���<��<���<���<s��<��<�	�<��<U)�<2�<�4�<2�<U)�<��<�	�<��<s��<���<���<��<���<'��<`   `   ]��<А�<��<���<'��<m��<���<��<p �<M5�<�E�<�O�<)S�<�O�<�E�<M5�<p �<��<���<m��<'��<���<��<А�<`   `   u��<���<��<H��<��<���<���<K�<;2�<*J�<�\�<rh�<�l�<rh�<�\�<*J�<;2�<K�<���<���<��<H��<��<���<`   `   b��<���<.��<]��<���<��<���<: �<�>�<CY�<�m�<{�<��<{�<�m�<CY�<�>�<: �<���<��<���<]��<.��<���<`   `   J}�<v��<h��<`��<���<r��<� �<P$�<CE�<�a�<x�<ޅ�<Ҋ�<ޅ�<x�<�a�<CE�<P$�<� �<r��<���<_��<h��<v��<`   `   �r�<Zw�<2��<���<��<@��</��<f"�<\E�<0c�<�z�<p��<���<p��<�z�<0c�<\E�<f"�</��<@��<��<���<2��<Zw�<`   `   Ff�<�j�<5y�<���<���<���<@��<o�<�?�<�]�<ov�<���<���<���<ov�<�]�<�?�<o�<@��<���<���<���<5y�<�j�<`   `   JX�<�\�<�j�<��<���<���<���<g�<�3�<mR�<	k�<�z�<��<�z�<	k�<mR�<�3�<g�<���<���<���<��<�j�<�\�<`   `   nI�<!N�<1\�<�r�<Y��<���<��<v��<	#�<.B�<1Z�<Vi�<�n�<Vi�<1Z�<.B�<	#�<v��<��<���<Y��<�r�<1\�<!N�<`   `   �:�<o?�<jM�<:c�<��<���<���<o��<$�<�-�<E�<mS�<�X�<mS�<E�<�-�<$�<o��<���<���<��<:c�<jM�<o?�<`   `   �-�<�1�<O?�<fT�<�o�<���<y��<`��<���<��<J,�<b:�<<?�<b:�<J,�<��<���<`��<y��<���<�o�<fT�<O?�<�1�<`   `   #�<%'�<�3�<�G�<ua�<��<��<q��<���<���<��<U�<�#�<U�<��<���<���<q��<��<��<ua�<�G�<�3�<%'�<`   `   ��<��<N+�<�=�<{U�<dq�<��<M��<]��<p��<i��<��<��<��<i��<p��<]��<M��<��<dq�<{U�<�=�<N+�<��<`   `   A?�<�B�<J�<V�<Ff�<�x�<���<���<��<���<��<J��<Q��<J��<��<���<��<���<���<�x�<Ff�<V�<J�<�B�<`   `   �A�<uD�<�J�</U�<5c�<�s�<I��<ۖ�<ݧ�<7��<H��<���<���<���<H��<7��<ݧ�<ۖ�<I��<�s�<5c�</U�<�J�<uD�<`   `   fH�<.J�<�O�< X�<%d�<�q�<���<���<���<���<��<f��<���<f��<��<���<���<���<���<�q�<%d�< X�<�O�<.J�<`   `   �R�<NT�<�X�<�_�<ki�<�s�<t�<X��<���<��<N��<a��<B��<a��<N��<��<���<X��<t�<�s�<ki�<�_�<�X�<NT�<`   `   �b�<Vc�<�f�<ok�<r�<�y�<���<���<���<[��<מ�<���<���<���<מ�<[��<���<���<���<�y�<r�<ok�<�f�<Vc�<`   `   v�<v�<�w�<�z�<�~�<;��<��<K��< ��<��<͙�<��< ��<��<͙�<��< ��<K��<��<;��<�~�<�z�<�w�<v�<`   `   Ό�<z��<
��<ލ�<���<��<2��<֒�<��<x��<��<���<ڗ�<���<��<x��<��<֒�<2��<��<���<ލ�<
��<z��<`   `   T��<˥�<���<T��<��<+��<��<���<���<���<���<r��<���<r��<���<���<���<���<��<+��<��<T��<���<˥�<`   `   ���<���</��<N��<b��<#��<>��<&��<?��<r��<ȗ�<���<@��<���<ȗ�<r��<?��<&��<>��<#��<b��<N��</��<���<`   `   :��<���<��<&��<���<���<)��<��<���<b��<��<���<v��<���<��<b��<���<��<)��<���<���<&��<��<���<`   `   j��<���<���<���<Y��<���<��<���<���<t��<v��<��<֕�<��<v��<t��<���<���<��<���<Y��<���<���<���<`   `   a�<��<�	�<^��< ��<���<���<+��<A��<Ч�<Ǟ�<��<���<��<Ǟ�<Ч�<A��<+��<���<���< ��<^��<�	�<��<`   `   �(�<�%�<D�<D�<��<��<��<(��<��<��<e��<z��<֕�<z��<e��<��<��<(��<��<��<��<D�<D�<�%�<`   `   /;�<
8�<�/�<�!�<��<���<���<Y��<���<���<W��<i��<���<i��<W��<���<���<Y��<���<���<��<�!�<�/�<
8�<`   `   �H�<`E�<$<�<-�<�<�<}��<���<���<F��<
��< ��<(��< ��<
��<F��<���<���<}��<�<�<-�<$<�<`E�<`   `   Q�<M�<+C�<>3�<��<��<��<���<Ѻ�<���<I��<S��<2��<S��<I��<���<Ѻ�<���<��<��<��<>3�<+C�<M�<`   `   T�<�O�<LE�<#4�<��<��<r��<���<;��<ޟ�<��<̅�<N��<̅�<��<ޟ�<;��<���<r��<��<��<#4�<LE�<�O�<`   `   �P�<%M�<MB�<�0�<��<4��<��<a��<���<���<��<z|�<�x�<z|�<��<���<���<a��<��<4��<��<�0�<MB�<%M�<`   `   aH�<�D�<:�<�(�<\�<*��<���<��<D��< ��<�|�<r�<Vn�<r�<�|�< ��<D��<��<���<*��<\�<�(�<:�<�D�<`   `   �<�<�8�<V-�<��<��</��<d��<U��<���<N��<�q�<)g�<rc�<)g�<�q�<N��<���<U��<d��</��<��<��<V-�<�8�<`   `   �,�<�(�<��<{�<���<Q��<��<̥�<8��<�v�<pf�<�[�<=X�<�[�<pf�<�v�<8��<̥�<��<Q��<���<{�<��<�(�<`   `   [�<��<��<O��<���<��<���<ј�<���<�k�<�[�<�Q�<�N�<�Q�<�[�<�k�<���<ј�<���<��<���<O��<��<��<`   `   G�<��<���<���<���<���<ݤ�<��<�u�<2b�<S�<@J�<bG�<@J�<S�<2b�<�u�<��<ݤ�<���<���<���<���<��<`   `   5��<���<���<��<5��<��<e��<#��<xl�<tZ�<�L�<�D�<�A�<�D�<�L�<tZ�<xl�<#��<e��<��<5��<��<���<���<`   `   Q��<J��<��<���<��<���<���<�x�<Ff�<V�<J�<�B�<A?�<�B�<J�<V�<Ff�<�x�<���<���<��<���<��<J��<`   `   ���<���<H��<7��<ݧ�<ۖ�<I��<�s�<5c�</U�<�J�<uD�<�A�<uD�<�J�</U�<5c�<�s�<I��<ۖ�<ݧ�<7��<H��<���<`   `   ���<f��<��<���<���<���<���<�q�<%d�< X�<�O�<.J�<fH�<.J�<�O�< X�<%d�<�q�<���<���<���<���<��<f��<`   `   B��<a��<N��<��<���<X��<t�<�s�<ki�<�_�<�X�<NT�<�R�<NT�<�X�<�_�<ki�<�s�<t�<X��<���<��<N��<a��<`   `   ���<���<מ�<[��<���<���<���<�y�<r�<ok�<�f�<Vc�<�b�<Vc�<�f�<ok�<r�<�y�<���<���<���<[��<מ�<���<`   `    ��<��<͙�<��< ��<K��<��<;��<�~�<�z�<�w�<v�<v�<v�<�w�<�z�<�~�<;��<��<K��< ��<��<͙�<��<`   `   ڗ�<���<��<x��<��<֒�<2��<��<���<ލ�<
��<z��<Ό�<z��<
��<ލ�<���<��<2��<֒�<��<x��<��<���<`   `   ���<r��<���<���<���<���<��<+��<��<T��<���<˥�<T��<˥�<���<T��<��<+��<��<���<���<���<���<r��<`   `   @��<���<ȗ�<r��<?��<&��<>��<#��<b��<N��</��<���<���<���</��<N��<b��<#��<>��<&��<?��<r��<ȗ�<���<`   `   v��<���<��<b��<���<��<)��<���<���<&��<��<���<:��<���<��<&��<���<���<)��<��<���<b��<��<���<`   `   ֕�<��<v��<t��<���<���<��<���<Y��<���<���<���<j��<���<���<���<Y��<���<��<���<���<t��<v��<��<`   `   ���<��<Ǟ�<Ч�<A��<+��<���<���< ��<^��<�	�<��<a�<��<�	�<^��< ��<���<���<+��<A��<Ч�<Ǟ�<��<`   `   ֕�<z��<e��<��<��<(��<��<��<��<D�<D�<�%�<�(�<�%�<D�<D�<��<��<��<(��<��<��<e��<z��<`   `   ���<i��<W��<���<���<Y��<���<���<��<�!�<�/�<
8�</;�<
8�<�/�<�!�<��<���<���<Y��<���<���<W��<i��<`   `   (��< ��<
��<F��<���<���<}��<�<�<-�<$<�<`E�<�H�<`E�<$<�<-�<�<�<}��<���<���<F��<
��< ��<`   `   2��<S��<I��<���<Ѻ�<���<��<��<��<>3�<+C�<M�<Q�<M�<+C�<>3�<��<��<��<���<Ѻ�<���<I��<S��<`   `   N��<̅�<��<ޟ�<;��<���<r��<��<��<#4�<LE�<�O�<T�<�O�<LE�<#4�<��<��<r��<���<;��<ޟ�<��<̅�<`   `   �x�<z|�<��<���<���<a��<��<4��<��<�0�<MB�<%M�<�P�<%M�<MB�<�0�<��<4��<��<a��<���<���<��<z|�<`   `   Vn�<r�<�|�< ��<D��<��<���<*��<\�<�(�<:�<�D�<aH�<�D�<:�<�(�<\�<*��<���<��<D��< ��<�|�<r�<`   `   rc�<)g�<�q�<N��<���<U��<d��</��<��<��<V-�<�8�<�<�<�8�<V-�<��<��</��<d��<U��<���<N��<�q�<)g�<`   `   =X�<�[�<pf�<�v�<8��<̥�<��<Q��<���<{�<��<�(�<�,�<�(�<��<{�<���<Q��<��<̥�<8��<�v�<pf�<�[�<`   `   �N�<�Q�<�[�<�k�<���<ј�<���<��<���<O��<��<��<[�<��<��<O��<���<��<���<ј�<���<�k�<�[�<�Q�<`   `   bG�<@J�<S�<2b�<�u�<��<ݤ�<���<���<���<���<��<G�<��<���<���<���<���<ݤ�<��<�u�<2b�<S�<@J�<`   `   �A�<�D�<�L�<tZ�<xl�<#��<e��<��<5��<��<���<���<5��<���<���<��<5��<��<e��<#��<xl�<tZ�<�L�<�D�<`   `   �[�<u]�<4c�<�l�<tx�<A��<��<��<D��<ݾ�<���<���<���<���<���<ݾ�<D��<��<��<A��<tx�<�l�<4c�<u]�<`   `   @]�<q^�<�c�<*l�<,v�<��<[��<���<��<���<8��<��<���<��<8��<���<��<���<[��<��<,v�<*l�<�c�<q^�<`   `   �a�<3c�<�g�<�n�<�v�<2��<.��<ږ�<��<`��<d��<h��<]��<h��<d��<`��<��<ږ�<.��<2��<�v�<�n�<�g�<3c�<`   `   �i�<Kk�<�n�<�s�<$z�<R��<Y��<��<��<���<���<��<ʭ�<��<���<���<��<��<Y��<R��<$z�<�s�<�n�<Kk�<`   `   @u�<Nv�<�x�<,|�<2��<܆�<+��<:��<>��<���</��<Τ�<��<Τ�</��<���<>��<:��<+��<܆�<2��<,|�<�x�<Nv�<`   `   ���<R��<���<���<Ŋ�<��<���<���<���<)��<��<���<u��<���<��<)��<���<���<���<��<Ŋ�<���<���<R��<`   `   ���<��<4��<Q��<4��<��<b��<Y��<���<ɛ�<��<���<1��<���<��<ɛ�<���<Y��<b��<��<4��<Q��<4��<��<`   `   ���<���<���<���<���<_��<��<���<��<���<���<W��<@��<W��<���<���<��<���<��<_��<���<���<���<���<`   `   ߻�<Z��<���<��<̳�<���<���<Ѧ�<���<���<՜�<���<z��<���<՜�<���<���<Ѧ�<���<���<̳�<��<���<Z��<`   `   ���<���<��<��<`��<��<=��<I��<��<���<���<@��<��<@��<���<���<��<I��<=��<��<`��<��<��<���<`   `   ���<���<"��<���<���<p��<���<��<���<���<e��<˜�<���<˜�<e��<���<���<��<���<p��<���<���<"��<���<`   `   ���<���<a��<��<,��<K��<��<���<���<U��<á�<G��<	��<G��<á�<U��<���<���<��<K��<,��<��<a��<���<`   `   a�<R�<� �<��<\��<?��<���<���<��<ت�<���<~��<��<~��<���<ت�<��<���<���<?��<\��<��<� �<R�<`   `   ��<��<��<]�<���<Z��<1��<c��<\��<ӫ�<���<h��<|��<h��<���<ӫ�<\��<c��<1��<Z��<���<]�<��<��<`   `   ��<��<|�<=�<G��<q��<���<]��<���<ܪ�<s��<z��<O��<z��<s��<ܪ�<���<]��<���<q��<G��<=�<|�<��<`   `   T&�<�#�<�<�<� �<���<g��<>��<ٶ�<Χ�<a��<G��<��<G��<a��<Χ�<ٶ�<>��<g��<���<� �<�<�<�#�<`   `   W(�<�%�<��<R�<� �<���<���<-��<���<���<+��<���<j��<���<+��<���<���<-��<���<���<� �<R�<��<�%�<`   `   G&�<#�<��<�<��<
��<j��<b��<֭�<:��<���<J��<k��<J��<���<:��<֭�<b��<j��<
��<��<�<��<#�<`   `   � �<��<��<��<���<s��<���<U��<��<=��<���<g��<V~�<g��<���<=��<��<U��<���<s��<���<��<��<��<`   `   ��<x�<"�<���<-��<���<���<ư�<���<��<���<�x�<v�<�x�<���<��<���<ư�<���<���<-��<���<"�<x�<`   `   �
�<{�<^ �<���<]��<(��<���<h��<��<̈́�<�x�<q�<�n�<q�<�x�<̈́�<��<h��<���<(��<]��<���<^ �<{�<`   `   ���<���<��<��<q��<���<6��<���<���<m|�<q�<�i�<g�<�i�<q�<m|�<���<���<6��<���<q��<��<��<���<`   `   ���<��<���<��<V��<"��<ܦ�<���<���<u�<@j�<$c�<�`�<$c�<@j�<u�<���<���<ܦ�<"��<V��<��<���<��<`   `   3��<	��<]��<5��< ��<Z��< ��<���<?}�<�o�<�e�<_�<�\�<_�<�e�<�o�<?}�<���< ��<Z��< ��<5��<]��<	��<`   `   ���<���<���<ܾ�<D��<��<��<A��<tx�<�l�<4c�<u]�<�[�<u]�<4c�<�l�<tx�<A��<��<��<D��<ݾ�<���<���<`   `   ���<��<8��<���<��<���<[��<��<,v�<*l�<�c�<q^�<@]�<q^�<�c�<*l�<,v�<��<[��<���<��<���<8��<��<`   `   ]��<h��<d��<`��<��<ږ�<.��<2��<�v�<�n�<�g�<3c�<�a�<3c�<�g�<�n�<�v�<2��<.��<ږ�<��<`��<d��<h��<`   `   ʭ�<��<���<���<��<��<Y��<R��<$z�<�s�<�n�<Kk�<�i�<Kk�<�n�<�s�<$z�<R��<Y��<��<��<���<���<��<`   `   ��<Τ�</��<���<>��<9��<+��<܆�<2��<,|�<�x�<Nv�<@u�<Nv�<�x�<,|�<2��<܆�<+��<9��<>��<���</��<Τ�<`   `   u��<���<��<)��<���<���<���<��<Ŋ�<���<���<R��<���<R��<���<���<Ŋ�<��<���<���<���<)��<��<���<`   `   1��<���<��<ɛ�<���<Y��<b��<��<4��<Q��<4��<��<���<��<4��<Q��<4��<��<b��<Y��<���<ɛ�<��<���<`   `   @��<W��<���<���<��<���<��<_��<���<���<���<���<���<���<���<���<���<_��<��<���<��<���<���<W��<`   `   z��<���<՜�<���<���<Ѧ�<���<���<̳�<��<���<Z��<߻�<Z��<���<��<̳�<���<���<Ѧ�<���<���<՜�<���<`   `   ��<@��<���<���<��<I��<=��<��<`��<��<��<���<���<���<��<��<`��<��<=��<I��<��<���<���<@��<`   `   ���<˜�<e��<���<���<��<���<p��<���<���<"��<���<���<���<"��<���<���<p��<���<��<���<���<e��<˜�<`   `   	��<G��<á�<U��<���<���<��<K��<,��<��<a��<���<���<���<a��<��<,��<K��<��<���<���<U��<á�<G��<`   `   ��<~��<���<ت�<��<���<���<?��<\��<��<� �<R�<a�<R�<� �<��<\��<?��<���<���<��<ت�<���<~��<`   `   |��<h��<���<ӫ�<\��<c��<1��<Z��<���<]�<��<��<��<��<��<]�<���<Z��<1��<c��<\��<ӫ�<���<h��<`   `   O��<z��<s��<ܪ�<���<]��<���<q��<G��<=�<|�<��<��<��<|�<=�<G��<q��<���<]��<���<ܪ�<s��<z��<`   `   ��<G��<a��<Χ�<ٶ�<>��<g��<���<� �<�<�<�#�<T&�<�#�<�<�<� �<���<g��<>��<ٶ�<Χ�<a��<G��<`   `   j��<���<+��<���<���<-��<���<���<� �<R�<��<�%�<W(�<�%�<��<R�<� �<���<���<-��<���<���<+��<���<`   `   l��<J��<���<:��<֭�<b��<j��<
��<��<�<��<#�<G&�<#�<��<�<��<
��<j��<b��<֭�<:��<���<J��<`   `   V~�<g��<���<=��<��<U��<���<s��<���<��<��<��<� �<��<��<��<���<s��<���<U��<��<=��<���<g��<`   `   v�<�x�<���<��<���<ư�<���<���<-��<���<"�<x�<��<x�<"�<���<-��<���<���<ư�<���<��<���<�x�<`   `   �n�<q�<�x�<̈́�<��<h��<���<(��<]��<���<^ �<{�<�
�<{�<^ �<���<]��<(��<���<h��<��<̈́�<�x�<q�<`   `   g�<�i�<q�<m|�<���<���<6��<���<q��<��<��<���<���<���<��<��<q��<���<6��<���<���<m|�<q�<�i�<`   `   �`�<$c�<@j�<u�<���<���<ܦ�<"��<V��<��<���<��<���<��<���<��<V��<"��<ܦ�<���<���<u�<@j�<$c�<`   `   �\�<_�<�e�<�o�<?}�<���< ��<[��< ��<5��<]��<	��<3��<	��<]��<5��< ��<Z��< ��<���<?}�<�o�<�e�<_�<`   `   8p�<rq�<�u�<|�<���<��<ښ�<���<���<���<���<��<���<��<���<���<���<���<ښ�<��<���<|�<�u�<rq�<`   `   q�<Ur�<�u�<�{�<5��<ތ�<y��<a��<���<u��<���<"��<&��<"��<���<u��<���<a��<y��<ތ�<5��<�{�<�u�<Ur�<`   `   wt�<�u�<x�<�}�<��<���<���<��<���<\��<���<Y��<A��<Y��<���<\��<���<��<���<���<��<�}�<x�<�u�<`   `   �z�<{�<�}�<���<���<���<��<˙�<ğ�<��<H��<d��<���<d��<H��<��<ğ�<˙�<��<���<���<���<�}�<{�<`   `   ��<���<��<��<���<܏�<v��<t��<���<*��<���<<��<��<<��<���<*��<���<t��<v��<܏�<���<��<��<���<`   `   ���<%��<!��<	��<��<���<���<ך�<'��<F��<K��<\��<���<\��<K��<F��<'��<ך�<���<���<��<	��<!��<%��<`   `   O��<���<ך�<&��<���<+��<&��<���<X��<5��<ҟ�<0��<ٟ�<0��<ҟ�<5��<X��<���<&��<+��<���<&��<ך�<���<`   `   ���<X��<���<���<ݥ�<���<A��<���<��<2��<���<z��<���<z��<���<2��<��<���<A��<���<ݥ�<���<���<X��<`   `   ���<��<���<���<��<ϭ�<���<���<���<��<A��<��<4��<��<A��<��<���<���<���<ϭ�<��<���<���<��<`   `   ���<���<��<��<p��<���<���<D��<p��<~��<;��<U��<ߞ�<U��<;��<~��<p��<D��<���<���<p��<��<��<���<`   `   ���<���<���<���<���<(��<���<ײ�<j��<%��<¢�<A��<��<A��<¢�<%��<j��<ײ�<���<(��<���<���<���<���<`   `   n��<n��<���<S��<L��<���<1��<Ѹ�<p��<V��<1��<���<��<���<1��<V��<p��<Ѹ�<1��<���<L��<S��<���<n��<`   `   ���<���<;��<���<$��<?��<��<��<���<���<ۤ�<���<,��<���<ۤ�<���<���<��<��<?��<$��<���<;��<���<`   `   ���<V��<o��<A��<���<I��<>��<w��<״�<���<L��<~��<%��<~��<L��<���<״�<w��<>��<I��<���<A��<o��<V��<`   `   �<���<���<��<���<6��<2��<+��<H��<���<���<���<8��<���<���<���<H��<+��<2��<6��<���<��<���<���<`   `   k�<�<%��<K��<��<���<��<���<���<r��<C��<��<��<��<C��<r��<���<���<��<���<��<K��<%��<�<`   `   ~�<%�<o��<)��<7��<��<���<���<��<b��<o��<���<o��<���<o��<b��<��<���<���<��<7��<)��<o��<%�<`   `   ��<��<���<1��<���<��<���<��<���<���<F��<D��<N��<D��<F��<���<���<��<���<��<���<1��<���<��<`   `   }�<L��<B��<���<��<Q��<���<���<���<#��<���<���<Չ�<���<���<#��<���<���<���<Q��<��<���<B��<L��<`   `   ��<A��<���<���<���<��<q��<R��<1��<B��<���<c��<���<c��<���<B��<1��<R��<q��<��<���<���<���<A��<`   `   ���<���<��<y��<&��<;��<,��<%��<r��<g��<��<7�<�}�<7�<��<g��<r��<%��<,��<;��<&��<y��<��<���<`   `   ���<���<���<��<)��<���<���<��<���<-��<n�<�y�<x�<�y�<n�<-��<���<��<���<���<)��<��<���<���<`   `   ���<���<���<���<Z��<X��<��<L��<���<���<�z�<vu�<�s�<vu�<�z�<���<���<L��<��<X��<Z��<���<���<���<`   `   b��<���<!��<^��<��<#��<���<���<���<�~�<9w�<�r�<Dq�<�r�<9w�<�~�<���<���<���<#��<��<^��<!��<���<`   `   ���<��<���<���<���<���<ښ�<��<���<|�<�u�<rq�<8p�<rq�<�u�<|�<���<��<ښ�<���<���<���<���<��<`   `   &��<"��<���<u��<���<a��<y��<ތ�<5��<�{�<�u�<Ur�<q�<Ur�<�u�<�{�<5��<ތ�<y��<a��<���<u��<���<"��<`   `   A��<Y��<���<\��<���<��<���<���<��<�}�<x�<�u�<wt�<�u�<x�<�}�<��<���<���<��<���<\��<���<Y��<`   `   ���<d��<H��<��<ğ�<˙�<��<���<���<���<�}�<{�<�z�<{�<�}�<���<���<���<��<˙�<ğ�<��<H��<d��<`   `   ��<<��<���<*��<���<t��<v��<܏�<���<��<��<���<��<���<��<��<���<܏�<v��<t��<���<*��<���<<��<`   `   ���<\��<K��<F��<'��<ך�<���<���<��<	��<!��<%��<���<%��<!��<	��<��<���<���<ך�<'��<F��<K��<\��<`   `   ٟ�<0��<ҟ�<5��<X��<���<&��<+��<���<&��<ך�<���<O��<���<ך�<&��<���<+��<&��<���<X��<5��<ҟ�<0��<`   `   ���<z��<���<2��<��<���<A��<���<ݥ�<���<���<X��<���<X��<���<���<ݥ�<���<A��<���<��<2��<���<z��<`   `   4��<��<A��<��<���<���<���<ϭ�<��<���<���<��<���<��<���<���<��<ϭ�<���<���<���<��<A��<��<`   `   ߞ�<U��<;��<~��<p��<D��<���<���<p��<��<��<���<���<���<��<��<p��<���<���<D��<p��<~��<;��<U��<`   `   ��<A��<¢�<%��<j��<ײ�<���<(��<���<���<���<���<���<���<���<���<���<(��<���<ײ�<j��<%��<¢�<A��<`   `   ��<���<1��<V��<p��<Ѹ�<1��<���<L��<S��<���<n��<n��<n��<���<S��<L��<���<1��<Ѹ�<p��<V��<1��<���<`   `   ,��<���<ۤ�<���<���<��<��<?��<$��<���<;��<���<���<���<;��<���<$��<?��<��<��<���<���<ۤ�<���<`   `   %��<~��<L��<���<״�<w��<>��<I��<���<A��<o��<V��<���<V��<o��<A��<���<I��<>��<w��<״�<���<L��<~��<`   `   8��<���<���<���<H��<+��<2��<6��<���<��<���<���<�<���<���<��<���<6��<2��<+��<H��<���<���<���<`   `   ��<��<C��<r��<���<���<��<���<��<K��<%��<�<k�<�<%��<K��<��<���<��<���<���<r��<C��<��<`   `   o��<���<o��<b��<��<���<���<��<7��<)��<o��<%�<~�<%�<o��<)��<7��<��<���<���<��<b��<o��<���<`   `   N��<D��<F��<���<���<��<���<��<���<1��<���<��<��<��<���<1��<���<��<���<��<���<���<F��<D��<`   `   Չ�<���<���<#��<���<���<���<Q��<��<���<B��<L��<}�<L��<B��<���<��<Q��<���<���<���<#��<���<���<`   `   ���<c��<���<B��<1��<R��<q��<��<���<���<���<A��<��<A��<���<���<���<��<q��<R��<1��<B��<���<c��<`   `   �}�<7�<��<g��<r��<%��<,��<;��<&��<y��<��<���<���<���<��<y��<&��<;��<,��<%��<r��<g��<��<7�<`   `   x�<�y�<n�<-��<���<��<���<���<)��<��<���<���<���<���<���<��<)��<���<���<��<���<-��<n�<�y�<`   `   �s�<vu�<�z�<���<���<L��<��<X��<Z��<���<���<���<���<���<���<���<Z��<X��<��<L��<���<���<�z�<vu�<`   `   Dq�<�r�<9w�<�~�<���<���<���<#��<��<^��<!��<���<b��<���<!��<^��<��<#��<���<���<���<�~�<9w�<�r�<`   `   f}�<�~�<���<ȇ�<b��<���<A��<M��<��<��<��<j��<���<j��<��<��<��<M��<A��<���<b��<ȇ�<���<�~�<`   `   ~�<;��<��<G��<;��<]��<ʚ�<��<��<��<Z��<I��<%��<I��<Z��<��<��<��<ʚ�<]��<;��<G��<��<;��<`   `   W��<���<���<i��<q��<���<ژ�<��<��<���<���<��<���<��<���<���<��<��<ژ�<���<q��<i��<���<���<`   `   ��<҆�<���<̋�<n��<$��<���<#��<���<l��<ͨ�<���<��<���<ͨ�<l��<���<#��<���<$��<n��<̋�<���<҆�<`   `   ��<���<j��<X��<���<���<���<�<e��<���<F��<j��<ۦ�<j��<F��<���<e��<�<���<���<���<X��<j��<���<`   `   ���<���<5��<V��<���<��<���<���<��<���<��<ţ�<*��<ţ�<��<���<��<���<���<��<���<V��<5��<���<`   `   ��<���<��<e��<���<F��<ȟ�<���<��<F��<���<��<���<��<���<F��<��<���<ȟ�<F��<���<e��<��<���<`   `   [��<���<���<(��< ��<���<���<u��<���<���<-��<
��<��<
��<-��<���<���<u��<���<���< ��<(��<���<���<`   `   ���<��<V��<y��<;��<o��<ک�<_��<_��<���<١�<��<C��<��<١�<���<_��<_��<ک�<o��<;��<y��<V��<��<`   `   Ͼ�< ��<���<\��<C��<���<���<��<i��<u��<��<g��<6��<g��<��<u��<i��<��<���<���<C��<\��<���< ��<`   `   ���<F��<���<���<v��<H��<��<.��<��<Ҧ�<A��<���<��<���<A��<Ҧ�<��<.��<��<H��<v��<���<���<F��<`   `   ���<���<���<f��<>��<���<g��<��<���<���< ��<m��<?��<m��< ��<���<���<��<g��<���<>��<f��<���<���<`   `   ���<��<��<C��<��<��<@��<9��<@��<��<t��<���<���<���<t��<��<@��<9��<@��<��<��<C��<��<��<`   `   ���<��<���<o��<���<A��<v��<;��<m��<o��<��<��<��<��<��<o��<m��<;��<v��<A��<���<o��<���<��<`   `   >��<v��<'��<Y��<���<���<5��<L��<���<��<���<{��<5��<{��<���<��<���<L��<5��<���<���<Y��<'��<v��<`   `   v��<���<���<���<���<��<���<E��<���<{��<A��<.��<���<.��<A��<{��<���<E��<���<��<���<���<���<���<`   `   ���<
��<T��<`��<���<���<���<ո�<R��<Υ�<<��<��<���<��<<��<Υ�<R��<ո�<���<���<���<`��<T��<
��<`   `   [��<���<v��<8��<S��<���<��<���<'��<J��<n��<F��<^��<F��<n��<J��<'��<���<��<���<S��<8��<v��<���<`   `   ��<>��<��<���<���<��<P��<F��<r��<M��<7��<֒�<ݑ�<֒�<7��<M��<r��<F��<P��<��<���<���<��<>��<`   `   ���<v��<���<���<���<-��<���<s��<s��<q��<���<|��<H��<|��<���<q��<s��<s��<���<-��<���<���<���<v��<`   `   E��<Z��<���<%��<��<|��<c��<��<b��<���<M��<:��<���<:��<M��<���<b��<��<c��<|��<��<%��<���<Z��<`   `   ���<���<u��<���<��<9��<���<ۢ�<0��<v��<��<���<:��<���<��<v��<0��<ۢ�<���<9��<��<���<u��<���<`   `   ���<���<���<_��<B��<��<���<^��<���<p��<5��<���<r��<���<5��<p��<���<^��<���<��<B��<_��<���<���<`   `   ��<���<���<��<���<��<���<��<���<K��<q��<��<�~�<��<q��<K��<���<��<���<��<���<��<���<���<`   `   ���<j��<��<��<��<M��<A��<���<b��<ȇ�<���<�~�<f}�<�~�<���<ȇ�<b��<���<A��<M��<��<��<��<j��<`   `   %��<I��<Z��<��<��<��<ʚ�<]��<;��<G��<��<;��<~�<;��<��<G��<;��<]��<ʚ�<��<��<��<Z��<I��<`   `   ���<��<���<���<��<��<ژ�<���<q��<i��<���<���<W��<���<���<i��<q��<���<ژ�<��<��<���<���<��<`   `   ��<���<ͨ�<l��<���<#��<���<$��<n��<̋�<���<҆�<��<҆�<���<̋�<n��<$��<���<#��<���<l��<ͨ�<���<`   `   ۦ�<j��<F��<���<e��<�<���<���<���<X��<j��<���<��<���<j��<X��<���<���<���<�<e��<���<F��<j��<`   `   *��<ţ�<��<���<��<���<���<��<���<V��<5��<���<���<���<5��<V��<���<��<���<���<��<���<��<ţ�<`   `   ���<��<���<F��<��<���<ȟ�<F��<���<e��<��<���<��<���<��<e��<���<F��<ȟ�<���<��<F��<���<��<`   `   ��<
��<-��<���<���<u��<���<���< ��<(��<���<���<[��<���<���<(��< ��<���<���<u��<���<���<-��<
��<`   `   C��<��<١�<���<_��<_��<ک�<o��<;��<y��<V��<��<���<��<V��<y��<;��<o��<ک�<_��<_��<���<١�<��<`   `   6��<g��<��<u��<i��<��<���<���<C��<\��<���< ��<Ͼ�< ��<���<\��<C��<���<���<��<i��<u��<��<g��<`   `   ��<���<A��<Ҧ�<��<.��<��<H��<v��<���<���<F��<���<F��<���<���<v��<H��<��<.��<��<Ҧ�<A��<���<`   `   ?��<m��< ��<���<���<��<g��<���<>��<f��<���<���<���<���<���<f��<>��<���<g��<��<���<���< ��<m��<`   `   ���<���<t��<��<@��<9��<@��<��<��<C��<��<��<���<��<��<C��<��<��<@��<9��<@��<��<t��<���<`   `   ��<��<��<o��<m��<;��<v��<A��<���<o��<���<��<���<��<���<o��<���<A��<v��<;��<m��<o��<��<��<`   `   5��<{��<���<��<���<L��<5��<���<���<Y��<'��<v��<>��<v��<'��<Y��<���<���<5��<L��<���<��<���<{��<`   `   ���<.��<A��<{��<���<E��<���<��<���<���<���<���<v��<���<���<���<���<��<���<E��<���<{��<A��<.��<`   `   ���<��<<��<Υ�<R��<ո�<���<���<���<`��<T��<
��<���<
��<T��<`��<���<���<���<ո�<R��<Υ�<<��<��<`   `   ^��<G��<n��<J��<'��<���<��<���<S��<8��<v��<���<[��<���<v��<8��<S��<���<��<���<'��<J��<n��<G��<`   `   ݑ�<֒�<7��<M��<r��<F��<P��<��<���<���<��<>��<��<>��<��<���<���<��<P��<F��<r��<M��<7��<֒�<`   `   H��<|��<���<q��<s��<s��<���<-��<���<���<���<v��<���<v��<���<���<���<-��<���<s��<s��<q��<���<|��<`   `   ���<:��<M��<���<b��<��<c��<|��<��<%��<���<Z��<E��<Z��<���<%��<��<|��<c��<��<b��<���<M��<:��<`   `   :��<���<��<v��<0��<ۢ�<���<9��<��<���<u��<���<���<���<u��<���<��<9��<���<ۢ�<0��<v��<��<���<`   `   r��<���<5��<p��<���<^��<���<��<B��<_��<���<���<���<���<���<_��<B��<��<���<^��<���<p��<5��<���<`   `   �~�<��<q��<K��<���<��<���<��<���<��<���<���<��<���<���<��<���<��<���<��<���<K��<q��<��<`   `   ߈�<?��<T��<���<G��<̙�<-��<p��<K��<b��<��<���<ӷ�<���<��<b��<K��<p��<-��<̙�<G��<���<T��<?��<`   `   T��<ǉ�<p��<���<^��<��<��<��<��<���<˯�<0��<,��<0��<˯�<���<��<��<��<��<^��<���<p��<ǉ�<`   `   ��<j��<���<ҏ�<]��<���<���<���<Τ�<���<7��<R��<s��<R��<7��<���<Τ�<���<���<���<]��<ҏ�<���<j��<`   `   ���<���<���<?��<���<ޗ�<���<C��<Ţ�<˥�<ǧ�<u��<
��<u��<ǧ�<˥�<Ţ�<C��<���<ޗ�<���<?��<���<���<`   `   ɒ�<#��<Z��<��<���<��<Ü�<E��<���<��<��<��<��<��<��<��<���<E��<Ü�<��<���<��<Z��<#��<`   `   ���<#��<�<g��<��<F��<t��<֟�<��<���<i��<��<���<��<i��<���<��<֟�<t��<F��<��<g��<�<#��<`   `   ��<��<��<C��<���<���<��<���<��<���<̢�<��<���<��<̢�<���<��<���<��<���<���<C��<��<��<`   `   ~��<U��<&��<��<H��<:��<���<l��<{��<���<���<;��<��<;��<���<���<{��<l��<���<:��<H��<��<&��<U��<`   `   ���<~��<���<���<k��<y��<���<���< ��<���<���<4��<$��<4��<���<���< ��<���<���<y��<k��<���<���<~��<`   `   ��<ڷ�<���<ڴ�<���<��<ج�<&��<{��</��<���<~��<(��<~��<���</��<{��<&��<ج�<��<���<ڴ�<���<ڷ�<`   `   B��<��<v��<��<��<V��<���<q��<,��<Ҧ�<t��<���<[��<���<t��<Ҧ�<,��<q��<���<V��<��<��<v��<��<`   `   ���<8��<e��<���<f��<&��<B��<د�<��<3��<ͤ�<C��<���<C��<ͤ�<3��<��<د�<B��<&��<f��<���<e��<8��<`   `   ���<���<���<9��<���<ݽ�<��<d��<j��<��<��<)��<���<)��<��<��<j��<d��<��<ݽ�<���<9��<���<���<`   `   q��<4��<���<h��<`��<��<���<Ĵ�<2��<��<Q��<Ƣ�<���<Ƣ�<Q��<��<2��<Ĵ�<���<��<`��<h��<���<4��<`   `   $��<���<p��<���<��<���<3��<b��<Y��<���<���<ˡ�<j��<ˡ�<���<���<Y��<b��<3��<���<��<���<p��<���<`   `   ���<Q��<���<���<���<z��<U��<��<��<���<���<��<���<��<���<���<��<��<U��<z��<���<���<���<Q��<`   `   ���<5��<��<'��<z��<���<»�<���<_��<��<���<���<Ϝ�<���<���<��<_��<���<»�<���<z��<'��<��<5��<`   `   s��<I��<2��<��<
��<j��<��<l��<��<���<���<5��<ę�<5��<���<���<��<l��<��<j��<
��<��<2��<I��<`   `   ��<��<���<���<z��<��<I��<���</��<<��<��<���<��<���<��<<��</��<���<I��<��<z��<���<���<��<`   `   p��<a��<"��<���<���<��<���<&��<���<Ϝ�<���<R��<��<R��<���<Ϝ�<���<&��<���<��<���<���<"��<a��<`   `   H��<r��<c��<P��<��<���<|��<X��<��<���<[��<��<ˏ�<��<[��<���<��<X��<|��<���<��<P��<c��<r��<`   `   ���<6��<5��<!��<��<R��<I��<���<,��<���<ɐ�<���<���<���<ɐ�<���<,��<���<I��<R��<��<!��<5��<6��<`   `   4��<y��<m��<}��<~��<���<��<��<���<���<f��<q��<\��<q��<f��<���<���<��<��<���<~��<}��<m��<y��<`   `   ���<7��<t��<K��<���<L��<l��<���<,��<���<���<��<��<��<���<���<,��<���<l��<L��<���<K��<t��<7��<`   `   ӷ�<���<��<b��<K��<p��<-��<̙�<G��<���<T��<?��<߈�<?��<T��<���<G��<̙�<-��<p��<K��<b��<��<���<`   `   ,��<0��<˯�<���<��<��<��<��<^��<���<p��<ǉ�<T��<ǉ�<p��<���<^��<��<��<��<��<���<˯�<0��<`   `   s��<R��<7��<���<Τ�<���<���<���<]��<ҏ�<���<j��<��<j��<���<ҏ�<]��<���<���<���<Τ�<���<7��<R��<`   `   
��<u��<ǧ�<˥�<Ţ�<C��<���<ޗ�<���<?��<���<���<���<���<���<?��<���<ޗ�<���<C��<Ţ�<˥�<ǧ�<u��<`   `   ��<��<��<��<���<E��<Ü�<��<���<��<Z��<#��<ɒ�<#��<Z��<��<���<��<Ü�<E��<���<��<��<��<`   `   ���<��<i��<���<��<֟�<t��<F��<��<g��<�<#��<���<#��<�<g��<��<F��<t��<֟�<��<���<i��<��<`   `   ���<��<̢�<���<��<���<��<���<���<C��<��<��<��<��<��<C��<���<���<��<���<��<���<̢�<��<`   `   ��<;��<���<���<{��<l��<���<:��<H��<��<&��<U��<~��<U��<&��<��<H��<:��<���<l��<{��<���<���<;��<`   `   $��<4��<���<���< ��<���<���<y��<k��<���<���<~��<���<~��<���<���<k��<y��<���<���< ��<���<���<4��<`   `   (��<~��<���</��<{��<&��<ج�<��<���<ڴ�<���<ڷ�<��<ڷ�<���<ڴ�<���<��<ج�<&��<{��</��<���<~��<`   `   [��<���<t��<Ҧ�<,��<q��<���<V��<��<��<v��<��<B��<��<v��<��<��<V��<���<q��<,��<Ҧ�<t��<���<`   `   ���<C��<ͤ�<3��<��<د�<B��<&��<f��<���<e��<8��<���<8��<e��<���<f��<&��<B��<د�<��<3��<ͤ�<C��<`   `   ���<)��<��<��<j��<d��<��<ݽ�<���<9��<���<���<���<���<���<9��<���<ݽ�<��<d��<j��<��<��<)��<`   `   ���<Ƣ�<Q��<��<2��<Ĵ�<���<��<`��<h��<���<4��<q��<4��<���<h��<`��<��<���<Ĵ�<2��<��<Q��<Ƣ�<`   `   j��<ˡ�<���<���<Y��<b��<3��<���<��<���<p��<���<$��<���<p��<���<��<���<3��<b��<Y��<���<���<ˡ�<`   `   ���<��<���<���<��<��<U��<z��<���<���<���<Q��<���<Q��<���<���<���<z��<U��<��<��<���<���<��<`   `   Ϝ�<���<���<��<_��<���<»�<���<z��<'��<��<5��<���<5��<��<'��<z��<���<»�<���<_��<��<���<���<`   `   ę�<5��<���<���<��<l��<��<j��<
��<��<2��<I��<s��<I��<2��<��<
��<j��<��<l��<��<���<���<5��<`   `   ��<���<��<<��</��<���<I��<��<z��<���<���<��<��<��<���<���<z��<��<I��<���</��<<��<��<���<`   `   ��<R��<���<Ϝ�<���<&��<���<��<���<���<"��<a��<p��<a��<"��<���<���<��<���<&��<���<Ϝ�<���<R��<`   `   ˏ�<��<[��<���<��<X��<|��<���<��<P��<c��<r��<H��<r��<c��<P��<��<���<|��<X��<��<���<[��<��<`   `   ���<���<ɐ�<���<,��<���<I��<R��<��<!��<5��<6��<���<6��<5��<!��<��<R��<I��<���<,��<���<ɐ�<���<`   `   \��<q��<f��<���<���<��<��<���<~��<}��<m��<y��<4��<y��<m��<}��<~��<���<��<��<���<���<f��<q��<`   `   ��<��<���<���<,��<���<l��<L��<���<K��<t��<7��<���<7��<t��<K��<���<L��<l��<���<,��<���<���<��<`   `   d��<|��<���<5��<ɗ�<+��<���<{��<���<J��<;��<a��<���<a��<;��<J��<���<{��<���<+��<ɗ�<5��<���<|��<`   `   v��<܏�<0��<Q��<P��<��<ڞ�<��<���<��<I��<:��<ܮ�<:��<I��<��<���<��<ڞ�<��<P��<Q��<0��<܏�<`   `   ���<a��<u��<-��<��<��<���<^��<���<���< ��<r��<��<r��< ��<���<���<^��<���<��<��<-��<u��<a��<`   `   ��<��<��<w��<��<(��<w��<���<Т�<��<���<���<��<���<���<��<Т�<���<w��<(��<��<w��<��<��<`   `   ,��<G��<���<��<��<*��<,��<���<ʡ�<Z��<ڤ�<q��<r��<q��<ڤ�<Z��<ʡ�<���<,��<*��<��<��<���<G��<`   `   3��<���<��<���<���<r��<ן�<��<͡�<���<���<ߣ�<���<ߣ�<���<���<͡�<��<ן�<r��<���<���<��<���<`   `   ���<Ҡ�<ʠ�<���<��<U��<ȡ�<���<D��<t��<���<���<â�<���<���<t��<D��<���<ȡ�<U��<��<���<ʠ�<Ҡ�<`   `   v��<o��<��<���<I��<��<���<���<i��<���<���<���<7��<���<���<���<i��<���<���<��<I��<���<��<o��<`   `   ���<���<ث�<��<��<ƨ�<���<+��<��<ݣ�<��<a��<��<a��<��<ݣ�<��<+��<���<ƨ�<��<��<ث�<���<`   `   ���<���<���<U��<���<m��<W��<P��<p��<���<F��<|��<S��<|��<F��<���<p��<P��<W��<m��<���<U��<���<���<`   `   ��<A��<?��<׵�<.��<e��<���<���<��<���<��<��<���<��<��<���<��<���<���<e��<.��<׵�<?��<A��<`   `   ��<ٽ�<R��<N��<L��<��<ʰ�<��<e��<���<���<O��<���<O��<���<���<e��<��<ʰ�<��<L��<N��<R��<ٽ�<`   `   |��<���<1��<L��<��<ڶ�<��<��<���<t��<פ�<@��<���<@��<פ�<t��<���<��<��<ڶ�<��<L��<1��<���<`   `   ��<���<N��<���<���<q��<���<1��<6��<���<���<٢�<��<٢�<���<���<6��<1��<���<q��<���<���<N��<���<`   `   ]��<���<���<��<N��<��<���<m��<[��<v��<��<"��<{��<"��<��<v��<[��<m��<���<��<N��<��<���<���<`   `   K��<���<F��<���<���<���<��<M��<��<���<��<��<���<��<��<���<��<M��<��<���<���<���<F��<���<`   `   ���<��<���<<��<-��<s��<��<���<é�<���<v��<)��<G��<)��<v��<���<é�<���<��<s��<-��<<��<���<��<`   `   &��<k��<���<��<��<��<B��<��<��<��<o��<��<��<��<o��<��<��<��<B��<��<��<��<���<k��<`   `   ���<���<���<^��<|��<C��<��<���<��<���<��<��<-��<��<��<���<��<���<��<C��<|��<^��<���<���<`   `   ���<��<���<���<׻�<���<���<L��<X��<R��<z��<y��<���<y��<z��<R��<X��<L��<���<���<׻�<���<���<��<`   `   @��<}��<��<��<��<{��<���<p��<���<���<Η�<���<��<���<Η�<���<���<p��<���<{��<��<��<��<}��<`   `   ���<j��<��<_��<���<\��<���<Z��<���<I��<l��<���<Q��<���<l��<I��<���<Z��<���<\��<���<_��<��<j��<`   `   ���<���<���<���<��<���<4��<���<T��<F��<��<���<���<���<��<F��<T��<���<4��<���<��<���<���<���<`   `   ���<0��<\��<a��<!��<M��</��<m��<u��<���<���<��<T��<��<���<���<u��<m��</��<M��<!��<a��<\��<0��<`   `   ���<a��<;��<J��<���<{��<���<+��<ɗ�<5��<���<|��<d��<|��<���<5��<ɗ�<+��<���<{��<���<J��<;��<a��<`   `   ܮ�<:��<I��<��<���<��<ڞ�<��<P��<Q��<0��<܏�<v��<܏�<0��<Q��<P��<��<ڞ�<��<���<��<I��<:��<`   `   ��<r��< ��<���<���<^��<���<��<��<-��<u��<a��<���<a��<u��<-��<��<��<���<^��<���<���< ��<r��<`   `   ��<���<���<��<Т�<���<w��<(��<��<w��<��<��<��<��<��<w��<��<(��<w��<���<Т�<��<���<���<`   `   r��<q��<ڤ�<Z��<ʡ�<���<,��<*��<��<��<���<G��<,��<G��<���<��<��<*��<,��<���<ʡ�<Z��<ڤ�<q��<`   `   ���<ߣ�<���<���<͡�<��<ן�<r��<���<���<��<���<3��<���<��<���<���<r��<ן�<��<͡�<���<���<ߣ�<`   `   â�<���<���<t��<D��<���<ȡ�<U��<��<���<ʠ�<Ҡ�<���<Ҡ�<ʠ�<���<��<U��<ȡ�<���<D��<t��<���<���<`   `   7��<���<���<���<i��<���<���<��<I��<���<��<o��<v��<o��<��<���<I��<��<���<���<i��<���<���<���<`   `   ��<a��<��<ݣ�<��<+��<���<ƨ�<��<��<ث�<���<���<���<ث�<��<��<ƨ�<���<+��<��<ݣ�<��<a��<`   `   S��<|��<F��<���<p��<P��<W��<m��<���<U��<���<���<���<���<���<U��<���<m��<W��<P��<p��<���<F��<|��<`   `   ���<��<��<���<��<���<���<e��<.��<׵�<?��<A��<��<A��<?��<׵�<.��<e��<���<���<��<���<��<��<`   `   ���<O��<���<���<e��<��<ʰ�<��<L��<N��<R��<ٽ�<��<ٽ�<R��<N��<L��<��<ʰ�<��<e��<���<���<O��<`   `   ���<@��<פ�<t��<���<��<��<ڶ�<��<L��<1��<���<|��<���<1��<L��<��<ڶ�<��<��<���<t��<פ�<@��<`   `   ��<٢�<���<���<6��<1��<���<q��<���<���<N��<���<��<���<N��<���<���<q��<���<1��<6��<���<���<٢�<`   `   {��<"��<��<v��<[��<m��<���<��<N��<��<���<���<]��<���<���<��<N��<��<���<m��<[��<v��<��<"��<`   `   ���<��<��<���<��<M��<��<���<���<���<F��<���<K��<���<F��<���<���<���<��<M��<��<���<��<��<`   `   G��<)��<v��<���<é�<���<��<s��<-��<<��<���<��<���<��<���<<��<-��<s��<��<���<é�<���<v��<)��<`   `   ��<��<o��<��<��<��<B��<��<��<��<���<k��<&��<k��<���<��<��<��<B��<��<��<��<o��<��<`   `   -��<��<��<���<��<���<��<C��<|��<^��<���<���<���<���<���<^��<|��<C��<��<���<��<���<��<��<`   `   ���<y��<z��<R��<X��<L��<���<���<׻�<���<���<��<���<��<���<���<׻�<���<���<L��<X��<R��<z��<y��<`   `    ��<���<Η�<���<���<p��<���<{��<��<��<��<}��<@��<}��<��<��<��<{��<���<p��<���<���<Η�<���<`   `   Q��<���<l��<I��<���<Z��<���<\��<���<_��<��<j��<���<j��<��<_��<���<\��<���<Z��<���<I��<l��<���<`   `   ���<���<��<F��<T��<���<4��<���<��<���<���<���<���<���<���<���<��<���<4��<���<T��<F��<��<���<`   `   T��<��<���<���<u��<m��</��<M��<!��<a��<\��<0��<���<0��<\��<a��<!��<M��</��<m��<u��<���<���<��<`   `   4��<��<���<ї�<���<؝�<4��<���<���<\��<��<~��<���<~��<��<\��<���<���<4��<؝�<���<ї�<���<��<`   `   ���<���<���<l��<��<���<���<Ң�<<��<ܧ�<���<{��<��<{��<���<ܧ�<<��<Ң�<���<���<��<l��<���<���<`   `   {��<���<k��<���<���<#��<���<���<���<���<`��<6��<���<6��<`��<���<���<���<���<#��<���<���<k��<���<`   `   ��<P��<N��<��<���<���<���<���<S��<���<��<���<(��<���<��<���<S��<���<���<���<���<��<N��<P��<`   `   ���<���<���<M��<9��<ȝ�<��<��<���<΢�<���<f��<o��<f��<���<΢�<���<��<��<ȝ�<9��<M��<���<���<`   `   ,��<'��<{��<��<Q��<-��<��<���<���<���<Т�<X��<^��<X��<Т�<���<���<���<��<-��<Q��<��<{��<'��<`   `   ܠ�<���<Ҡ�<X��<O��<���<���<���<]��<"��<��<u��<x��<u��<��<"��<]��<���<���<���<O��<X��<Ҡ�<���<`   `   ���<ݤ�<��<��<L��<��<O��<Ţ�<֢�<N��<��<&��<��<&��<��<N��<֢�<Ţ�<O��<��<L��<��<��<ݤ�<`   `   Y��<e��<,��<���<���<���<���<���<У�<��<b��<)��<+��<)��<b��<��<У�<���<���<���<���<���<,��<e��<`   `   ��<��<=��<&��<��<é�<L��<���<
��<��<��<H��<?��<H��<��<��<
��<���<L��<é�<��<&��<=��<��<`   `   ���<a��<���<"��<���<���<!��<S��<C��<���<���<o��<��<o��<���<���<C��<S��<!��<���<���<"��<���<a��<`   `   ���<|��<���<ճ�<ڱ�<3��<)��<��<e��<7��<̣�<x��<ҡ�<x��<̣�<7��<e��<��<)��<3��<ڱ�<ճ�<���<|��<`   `   H��<��<���<���<C��<���<D��<��<C��<¥�<٣�<���</��<���<٣�<¥�<C��<��<D��<���<C��<���<���<��<`   `   _��<Ƽ�<{��<M��<U��<Z��<���<���<ܨ�<��<���<���<F��<���<���<��<ܨ�<���<���<Z��<U��<M��<{��<Ƽ�<`   `   ���<��<q��<���<ҷ�<+��<���<^��<��<ҥ�<���<���<!��<���<���<ҥ�<��<^��<���<+��<ҷ�<���<q��<��<`   `   ��<h��<���<R��<���<���<���<_��<���<%��<���<Š�<���<Š�<���<%��<���<_��<���<���<���<R��<���<h��<`   `   #��<���<��<A��<���<ٴ�<��<���<���<&��<���<���<&��<���<���<&��<���<���<��<ٴ�<���<A��<��<���<`   `   ���<���<���<���<��<߳�<���<���<���<��<ڟ�<��<��<��<ڟ�<��<���<���<���<߳�<��<���<���<���<`   `   ���<��<��<N��<���<0��<���<��<��<_��<7��<��<���<��<7��<_��<��<��<���<0��<���<N��<��<��<`   `   ���<��<+��<u��<���<W��<���<��<���<>��<���<F��<���<F��<���<>��<���<��<���<W��<���<u��<+��<��<`   `   G��<m��<��<��<H��<��<;��<���<���<	��<���<���<w��<���<���<	��<���<���<;��<��<H��<��<��<m��<`   `   ��<��<��<4��<���<���<���<Т�<��<p��<Ø�<��<��<��<Ø�<p��<��<Т�<���<���<���<4��<��<��<`   `   ڴ�<��<���<��<���<
��<ʤ�<���<��<���<ߖ�<���<��<���<ߖ�<���<��<���<ʤ�<
��<���<��<���<��<`   `   ı�<0��<���<��<��<���<Ģ�<ɞ�<Z��<C��<���<���<O��<���<���<C��<Z��<ɞ�<Ģ�<���<��<��<���<0��<`   `   ���<~��<��<\��<���<���<4��<؝�<���<ї�<���<��<4��<��<���<ї�<���<؝�<4��<���<���<\��<��<~��<`   `   ��<{��<���<ܧ�<<��<Ң�<���<���<��<l��<���<���<���<���<���<l��<��<���<���<Ң�<<��<ܧ�<���<{��<`   `   ���<6��<`��<���<���<���<���<#��<���<���<k��<���<{��<���<k��<���<���<#��<���<���<���<���<`��<6��<`   `   (��<���<��<���<S��<���<���<���<���<��<N��<P��<��<P��<N��<��<���<���<���<���<S��<���<��<���<`   `   o��<f��<���<΢�<���<��<��<ȝ�<9��<M��<���<���<���<���<���<M��<9��<ȝ�<��<��<���<΢�<���<f��<`   `   ^��<X��<Т�<���<���<���<��<-��<Q��<��<{��<'��<,��<'��<{��<��<Q��<-��<��<���<���<���<Т�<X��<`   `   x��<u��<��<"��<]��<���<���<���<O��<X��<Ҡ�<���<ܠ�<���<Ҡ�<X��<O��<���<���<���<]��<"��<��<u��<`   `   ��<&��<��<N��<֢�<Ţ�<O��<��<L��<��<��<ݤ�<���<ݤ�<��<��<L��<��<O��<Ţ�<֢�<N��<��<&��<`   `   +��<)��<b��<��<У�<���<���<���<���<���<,��<e��<Y��<e��<,��<���<���<���<���<���<У�<��<b��<)��<`   `   ?��<H��<��<��<
��<���<L��<é�<��<&��<=��<��<��<��<=��<&��<��<é�<L��<���<
��<��<��<H��<`   `   ��<o��<���<���<C��<S��<!��<���<���<"��<���<a��<���<a��<���<"��<���<���<!��<S��<C��<���<���<o��<`   `   ҡ�<x��<̣�<7��<e��<��<)��<3��<ڱ�<ճ�<���<|��<���<|��<���<ճ�<ڱ�<3��<)��<��<e��<7��<̣�<x��<`   `   /��<���<٣�<¥�<C��<��<D��<���<C��<���<���<��<H��<��<���<���<C��<���<D��<��<C��<¥�<٣�<���<`   `   F��<���<���<��<ܨ�<���<���<Z��<U��<M��<{��<Ƽ�<_��<Ƽ�<{��<M��<U��<Z��<���<���<ܨ�<��<���<���<`   `   !��<���<���<ҥ�<��<^��<���<+��<ҷ�<���<q��<��<���<��<q��<���<ҷ�<+��<���<^��<��<ҥ�<���<���<`   `   ���<Š�<���<%��<���<_��<���<���<���<R��<���<h��<��<h��<���<R��<���<���<���<_��<���<%��<���<Š�<`   `   &��<���<���<&��<���<���<��<ٴ�<���<A��<��<���<#��<���<��<A��<���<ٴ�<��<���<���<&��<���<���<`   `   ��<��<ڟ�<��<���<���<���<߳�<��<���<���<���<���<���<���<���<��<߳�<���<���<���<��<ڟ�<��<`   `   ���<��<7��<_��<��<��<���<0��<���<N��<��<��<���<��<��<N��<���<0��<���<��<��<_��<7��<��<`   `   ���<F��<���<>��<���<��<���<W��<���<u��<+��<��<���<��<+��<u��<���<W��<���<��<���<>��<���<F��<`   `   w��<���<���<	��<���<���<;��<��<H��<��<��<m��<G��<m��<��<��<H��<��<;��<���<���<	��<���<���<`   `   ��<��<Ø�<p��<��<Т�<���<���<���<4��<��<��<��<��<��<4��<���<���<���<Т�<��<p��<Ø�<��<`   `   ��<���<ߖ�<���<��<���<ʤ�<
��<���<��<���<��<ڴ�<��<���<��<���<
��<ʤ�<���<��<���<ߖ�<���<`   `   O��<���<���<C��<Z��<ɞ�<Ģ�<���<��<��<���<0��<ı�<0��<���<��<��<���<Ģ�<ɞ�<Z��<C��<���<���<`   `   ̕�<��<��<���<o��<Ý�<W��<���<x��<y��<ר�<���<*��<���<ר�<y��<x��<���<W��<Ý�<o��<���<��<��<`   `   ���<6��<˗�<���<W��<L��<���<w��<���<j��<��<���<F��<���<��<j��<���<w��<���<L��<W��<���<˗�<6��<`   `   '��<+��<���<D��<���<՜�<Ԟ�<���<D��<���<��<¥�<��<¥�<��<���<D��<���<Ԟ�<՜�<���<D��<���<+��<`   `   ۘ�<2��<��<G��<���<0��<ߞ�<!��<ء�<��<���<��<6��<��<���<��<ء�<!��<ߞ�<0��<���<G��<��<2��<`   `   ��<��<g��<7��<Ӝ�<��<>��<��<R��<!��<d��<��<+��<��<d��<!��<R��<��<>��<��<Ӝ�<7��<g��<��<`   `   ���<u��<v��<��<���<��<���<C��<���<9��<���<ҡ�<��<ҡ�<���<9��<���<C��<���<��<���<��<v��<u��<`   `   ]��<]��<X��<T��<���<���<ߠ�<h��<֠�<B��<֡�<Z��<q��<Z��<֡�<B��<֠�<h��<ߠ�<���<���<T��<X��<]��<`   `   Σ�<���<L��<���<���<���<G��<���<���<���<ҡ�<-��<#��<-��<ҡ�<���<���<���<G��<���<���<���<L��<���<`   `   ��<���<Y��<��<{��<���<ϣ�<N��<{��<ڡ�<���<��<��<��<���<ڡ�<{��<N��<ϣ�<���<{��<��<Y��<���<`   `   s��<,��<���<��<��<���<̥�<v��<G��<^��<���<M��<��<M��<���<^��<G��<v��<̥�<���<��<��<���<,��<`   `   ���<v��<Ƭ�<��<D��<��<���<��<H��<��< ��<���<���<���< ��<��<H��<��<���<��<D��<��<Ƭ�<v��<`   `   b��<-��<���<d��<ì�<��<��<"��<7��<���<I��<���<��<���<I��<���<7��<"��<��<��<ì�<d��<���<-��<`   `   ���<��<��<���<��<���<A��<��<��<ޣ�<}��<���<[��<���<}��<ޣ�<��<��<A��<���<��<���<��<��<`   `   ��<]��<���<���<6��<׭�<J��<���<[��<���<���<w��<ɠ�<w��<���<���<[��<���<J��<׭�<6��<���<���<]��<`   `   ��<޶�<���<��<���<ۮ�<��<��<Q��<���<���<h��<���<h��<���<���<Q��<��<��<ۮ�<���<��<���<޶�<`   `   ���<˷�<���<���<%��<U��<
��<	��<���<.��<���<r��<
��<r��<���<.��<���<	��<
��<U��<%��<���<���<˷�<`   `   x��<���<���<���<��<��<p��<���<u��<���<���<g��<T��<g��<���<���<u��<���<p��<��<��<���<���<���<`   `   0��<���<���<���<z��<���<��<ç�<@��<z��<���<K��<-��<K��<���<z��<@��<ç�<��<���<z��<���<���<���<`   `   ;��<���<���<���<O��<r��<��<^��<٢�<J��<u��<ڜ�<���<ڜ�<u��<J��<٢�<^��<��<r��<O��<���<���<���<`   `   ��<E��<��<���<ڮ�<��<g��<��<��<���<��<���<���<���<��<���<��<��<g��<��<ڮ�<���<��<E��<`   `   ��<s��<��<��<b��<j��<¦�<���<o��<X��<|��<���<l��<���<|��<X��<o��<���<¦�<j��<b��<��<��<s��<`   `   x��<4��<���<��<_��<D��<��<���<���<��<U��<	��<`��<	��<U��<��<���<���<��<D��<_��<��<���<4��<`   `   ���<��<���<n��<U��<N��<���<t��<~��<��<��< ��<a��< ��<��<��<~��<t��<���<N��<U��<n��<���<��<`   `   ���<[��<��<M��<p��<G��<���<Ş�<1��<��<k��<���<ʖ�<���<k��<��<1��<Ş�<���<G��<p��<M��<��<[��<`   `   *��<���<ר�<x��<x��<���<W��<Ý�<o��<���<��<��<̕�<��<��<���<o��<Ý�<W��<���<x��<x��<ר�<���<`   `   F��<���<��<j��<���<w��<���<L��<W��<���<˗�<6��<���<6��<˗�<���<W��<L��<���<w��<���<j��<��<���<`   `   ��<¥�<��<���<D��<���<Ԟ�<՜�<���<D��<���<+��<'��<+��<���<D��<���<՜�<Ԟ�<���<D��<���<��<¥�<`   `   6��<��<���<��<ء�<!��<ߞ�<0��<���<G��<��<2��<ۘ�<2��<��<G��<���<0��<ߞ�<!��<ء�<��<���<��<`   `   +��<��<d��<!��<R��<��<>��<��<Ӝ�<7��<g��<��<��<��<g��<7��<Ӝ�<��<>��<��<R��<!��<d��<��<`   `   ��<ҡ�<���<9��<���<C��<���<��<���<��<v��<u��<���<u��<v��<��<���<��<���<C��<���<9��<���<ҡ�<`   `   q��<Z��<֡�<B��<֠�<h��<ߠ�<���<���<T��<X��<]��<]��<]��<X��<T��<���<���<ߠ�<h��<֠�<B��<֡�<Z��<`   `   #��<-��<ҡ�<���<���<���<G��<���<���<���<L��<���<Σ�<���<L��<���<���<���<G��<���<���<���<ҡ�<-��<`   `   ��<��<���<ڡ�<{��<N��<ϣ�<���<{��<��<Y��<���<��<���<Y��<��<{��<���<ϣ�<N��<{��<ڡ�<���<��<`   `   ��<M��<���<^��<G��<v��<̥�<���<��<��<���<,��<s��<,��<���<��<��<���<̥�<v��<G��<^��<���<M��<`   `   ���<���< ��<��<H��<��<���<��<D��<��<Ƭ�<v��<���<v��<Ƭ�<��<D��<��<���<��<H��<��< ��<���<`   `   ��<���<I��<���<7��<"��<��<��<ì�<d��<���<-��<b��<-��<���<d��<ì�<��<��<"��<7��<���<I��<���<`   `   [��<���<}��<ޣ�<��<��<A��<���<��<���<��<��<���<��<��<���<��<���<A��<��<��<ޣ�<}��<���<`   `   ɠ�<w��<���<���<[��<���<J��<׭�<6��<���<���<]��<��<]��<���<���<6��<׭�<J��<���<[��<���<���<w��<`   `   ���<h��<���<���<Q��<��<��<ۮ�<���<��<���<޶�<��<޶�<���<��<���<ۮ�<��<��<Q��<���<���<h��<`   `   
��<r��<���<.��<���<	��<
��<U��<%��<���<���<˷�<���<˷�<���<���<%��<U��<
��<	��<���<.��<���<r��<`   `   T��<g��<���<���<u��<���<p��<��<��<���<���<���<x��<���<���<���<��<��<p��<���<u��<���<���<g��<`   `   -��<K��<���<z��<@��<ç�<��<���<z��<���<���<���<0��<���<���<���<z��<���<��<ç�<@��<z��<���<K��<`   `   ���<ڜ�<u��<J��<٢�<^��<��<r��<O��<���<���<���<;��<���<���<���<O��<r��<��<^��<٢�<J��<u��<ڜ�<`   `   ���<���<��<���<��<��<g��<��<ڮ�<���<��<E��<��<E��<��<���<ڮ�<��<g��<��<��<���<��<���<`   `   l��<���<|��<X��<o��<���<¦�<j��<b��<��<��<s��<��<s��<��<��<b��<j��<¦�<���<o��<X��<|��<���<`   `   `��<	��<U��<��<���<���<��<D��<_��<��<���<4��<x��<4��<���<��<_��<D��<��<���<���<��<U��<	��<`   `   a��< ��<��<��<~��<t��<���<N��<U��<n��<���<��<���<��<���<n��<U��<N��<���<t��<~��<��<��< ��<`   `   ʖ�<���<k��<��<1��<Ş�<���<G��<p��<M��<��<[��<���<[��<��<M��<p��<G��<���<Ş�<1��<��<k��<���<`   `   ;��<���<)��<_��<���<���<���<j��<"��<o��<٥�<���<��<���<٥�<o��<"��<j��<���<���<���<_��<)��<���<`   `   j��<���<p��<8��<[��<9��<��<���<W��<;��<D��<��<9��<��<D��<;��<W��<���<��<9��<[��<8��<p��<���<`   `   ј�<n��<ҙ�<���<���<%��<s��<���<7��<��<��<A��<]��<A��<��<��<7��<���<s��<%��<���<���<ҙ�<n��<`   `   ��<e��<q��<��<��<���<��<��<!��<��<���<_��<e��<_��<���<��<!��<��<��<���<��<��<q��<e��<`   `   қ�<��<ћ�<:��<$��<���<~��<c��<��<_��<0��<���<���<���<0��<_��<��<c��<~��<���<$��<:��<ћ�<��<`   `   %��<u��<���<���<x��<���<���<ڟ�<���<1��<���<���<à�<���<���<1��<���<ڟ�<���<���<x��<���<���<u��<`   `   ��<d��<��<���<���<���<~��<��<���<U��<H��<1��<Ġ�<1��<H��<U��<���<��<~��<���<���<���<��<d��<`   `   ���<¡�<ݡ�<w��<w��<z��<���<���<[��<Z��<��<��<���<��<��<Z��<[��<���<���<z��<w��<w��<ݡ�<¡�<`   `   6��<��<ݣ�<���<E��<٢�<8��<���<F��<���<,��<B��<3��<B��<,��<���<F��<���<8��<٢�<E��<���<ݣ�<��<`   `   ���<���<\��<��<���<���<:��<n��<��<2��<���<���<���<���<���<2��<��<n��<:��<���<���<��<\��<���<`   `   2��<��<���< ��<��<��<ˤ�<d��<���<���<���<4��<͟�<4��<���<���<���<d��<ˤ�<��<��< ��<���<��<`   `   ���<a��<���<٩�<���<S��<��<9��<آ�<��<!��<V��<G��<V��<!��<��<آ�<9��<��<S��<���<٩�<���<a��<`   `   x��<S��<���<���<'��<���<	��<7��<a��</��<^��<c��<Y��<c��<^��</��<a��<7��<	��<���<'��<���<���<S��<`   `   ���<���<��<��<���<���<���<ե�<ѣ�<!��<��<��<��<��<��<!��<ѣ�<ե�<���<���<���<��<��<���<`   `   ɯ�<A��<6��<���<Q��<+��<���<ť�<ɣ�<9��<ߠ�<џ�<��<џ�<ߠ�<9��<ɣ�<ť�<���<+��<Q��<���<6��<A��<`   `   ��<���<���<S��<���<���<��<���<���<��<S��<?��<j��<?��<S��<��<���<���<��<���<���<S��<���<���<`   `   ±�<���<��<���<��<.��<���<|��<B��<���<���<���<b��<���<���<���<B��<|��<���<.��<��<���<��<���<`   `   S��<s��<h��<2��<E��<���<Z��<��<���<���<��<(��<R��<(��<��<���<���<��<Z��<���<E��<2��<h��<s��<`   `   ���<��<ʮ�<U��<���<��<P��<��<���<}��<!��<D��<X��<D��<!��<}��<���<��<P��<��<���<U��<ʮ�<��<`   `   ��<��<��<u��<i��<ۧ�<V��<͢�<Ҡ�<���<؜�<��<��<��<؜�<���<Ҡ�<͢�<V��<ۧ�<i��<u��<��<��<`   `   r��<p��<v��<��<��<���<[��<���<x��<���<ћ�<���<���<���<ћ�<���<x��<���<[��<���<��<��<v��<p��<`   `   X��<��<Ȫ�<���<v��<��<ۢ�<3��<��<���<��<Й�<��<Й�<��<���<��<3��<ۢ�<��<v��<���<Ȫ�<��<`   `   `��<&��<-��<��<8��<ڣ�<���<g��<K��<���<#��<!��<1��<!��<#��<���<K��<g��<���<ڣ�<8��<��<-��<&��<`   `   a��<-��<{��<;��<���<���<���<���<ɜ�<��<S��<���<���<���<S��<��<ɜ�<���<���<���<���<;��<{��<-��<`   `   ��<���<٥�<o��<"��<j��<���<���<���<_��<)��<���<;��<���<)��<_��<���<���<���<j��<"��<o��<٥�<���<`   `   9��<��<C��<;��<W��<���<��<9��<[��<8��<p��<���<j��<���<p��<8��<[��<9��<��<���<W��<;��<C��<��<`   `   ]��<A��<��<��<7��<���<s��<%��<���<���<ҙ�<n��<ј�<n��<ҙ�<���<���<%��<s��<���<7��<��<��<A��<`   `   e��<_��<���<��<!��<��<��<���<��<��<q��<e��<��<e��<q��<��<��<���<��<��<!��<��<���<_��<`   `   ���<���<0��<_��<��<c��<~��<���<$��<:��<ћ�<��<қ�<��<ћ�<:��<$��<���<~��<c��<��<_��<0��<���<`   `   à�<���<���<1��<���<ڟ�<���<���<x��<���<���<u��<%��<u��<���<���<x��<���<���<ڟ�<���<1��<���<���<`   `   Ġ�<1��<H��<U��<���<��<~��<���<���<���<��<d��<��<d��<��<���<���<���<~��<��<���<U��<H��<1��<`   `   ���<��<��<Z��<[��<���<���<z��<w��<w��<ݡ�<¡�<���<¡�<ݡ�<w��<w��<z��<���<���<[��<Z��<��<��<`   `   3��<B��<,��<���<F��<���<8��<٢�<E��<���<ݣ�<��<6��<��<ݣ�<���<E��<٢�<8��<���<F��<���<,��<B��<`   `   ���<���<���<2��<��<n��<:��<���<���<��<\��<���<���<���<\��<��<���<���<:��<n��<��<2��<���<���<`   `   ͟�<4��<���<���<���<d��<ˤ�<��<��< ��<���<��<2��<��<���< ��<��<��<ˤ�<d��<���<���<���<4��<`   `   G��<V��<!��<��<آ�<9��<��<S��<���<٩�<���<a��<���<a��<���<٩�<���<S��<��<9��<آ�<��<!��<V��<`   `   Y��<c��<^��</��<a��<7��<	��<���<'��<���<���<S��<x��<S��<���<���<'��<���<	��<7��<a��</��<^��<c��<`   `   ��<��<��<!��<ѣ�<ե�<���<���<���<��<��<���<���<���<��<��<���<���<���<ե�<ѣ�<!��<��<��<`   `   ��<џ�<ߠ�<9��<ɣ�<ť�<���<+��<Q��<���<6��<A��<ɯ�<A��<6��<���<Q��<+��<���<ť�<ɣ�<9��<ߠ�<џ�<`   `   j��<?��<S��<��<���<���<��<���<���<S��<���<���<��<���<���<S��<���<���<��<���<���<��<S��<?��<`   `   b��<���<���<���<B��<|��<���<.��<��<���<��<���<±�<���<��<���<��<.��<���<|��<B��<���<���<���<`   `   R��<(��<��<���<���<��<Z��<���<E��<2��<h��<s��<S��<s��<h��<2��<E��<���<Z��<��<���<���<��<(��<`   `   X��<D��<!��<}��<���<��<P��<��<���<U��<ʮ�<��<���<��<ʮ�<U��<���<��<P��<��<���<}��<!��<D��<`   `   ��<��<؜�<���<Ҡ�<͢�<V��<ۧ�<i��<u��<��<��<��<��<��<u��<i��<ۧ�<V��<͢�<Ҡ�<���<؜�<��<`   `   ���<���<ћ�<���<x��<���<[��<���<��<��<v��<p��<r��<p��<v��<��<��<���<[��<���<x��<���<ћ�<���<`   `   ��<Й�<��<���<��<4��<ۢ�<��<v��<���<Ȫ�<��<X��<��<Ȫ�<���<v��<��<ۢ�<4��<��<���<��<Й�<`   `   1��<!��<#��<���<K��<g��<���<ڣ�<8��<��<-��<&��<`��<&��<-��<��<8��<ڣ�<���<g��<K��<���<#��<!��<`   `   ���<���<S��<	��<ɜ�<���<���<���<���<;��<{��<-��<a��<-��<{��<;��<���<���<���<���<ɜ�<	��<S��<���<`   `   ���<)��<���<���<ޛ�<��<@��<��<Ơ�<��<(��<`��<���<`��<(��<��<Ơ�<��<@��<��<ޛ�<���<���<)��<`   `   L��<��<���<���<��<���<e��<̞�<��<��<��<%��<"��<%��<��<��<��<̞�<e��<���<��<���<���<��<`   `   \��<}��<$��<���<o��<���<j��<o��<^��<P��<���<k��<���<k��<���<P��<^��<o��<j��<���<o��<���<$��<}��<`   `   H��<j��<ך�<+��<��<���<���<x��<��<���<��<P��<���<P��<��<���<��<x��<���<���<��<+��<ך�<j��<`   `   ��<?��<��<4��<���<��<h��<��<���<��<a��<���<��<���<a��<��<���<��<h��<��<���<4��<��<?��<`   `   Ɯ�<���<Ɯ�<���<��<ם�<��<��<Ȟ�<��<��<F��<��<F��<��<��<Ȟ�<��<��<ם�<��<���<Ɯ�<���<`   `   ��<L��<��<;��<��<���<���<���<��<��<Ş�<��<Ӟ�<��<Ş�<��<��<���<���<���<��<;��<��<L��<`   `   /��<��<���<"��<���<\��<l��<��<��<���<͞�<˞�<���<˞�<͞�<���<��<��<l��<\��<���<"��<���<��<`   `   ��<���<���<Y��<��<���<s��<̟�<f��<.��<���<���<N��<���<���<.��<f��<̟�<s��<���<��<Y��<���<���<`   `   ˣ�<ƣ�<\��<���<V��<ء�<X��<���<ӟ�<G��<���<��<���<��<���<G��<ӟ�<���<X��<ء�<V��<���<\��<ƣ�<`   `   H��<\��<��<���<<��<4��<9��<~��<���<���<��<��<؞�<��<��<���<���<~��<9��<4��<<��<���<��<\��<`   `   G��<F��<̦�<��< ��<��<ʢ�<���<��<��<_��<���<���<���<_��<��<��<���<ʢ�<��< ��<��<̦�<F��<`   `   ���<���<	��<��<���<��<���<N��<f��<0��<p��<��<���<��<p��<0��<f��<N��<���<��<���<��<	��<���<`   `   ���<ѩ�<;��<]��<��<��<a��<Т�<���<T��<d��<���<-��<���<d��<T��<���<Т�<a��<��<��<]��<;��<ѩ�<`   `   C��<���<��<��<���<��<���<&��<���<^��<7��<���<���<���<7��<^��<���<&��<���<��<���<��<��<���<`   `   Z��<���<8��<z��<��<W��<���<.��<P��<���<��<m��<��<m��<��<���<P��<.��<���<W��<��<z��<8��<���<`   `   l��<��<ժ�<���<��<U��<���<���<���<t��<g��<9��<���<9��<g��<t��<���<���<���<U��<��<���<ժ�<��<`   `   ��<8��<���<���<ا�<���<��<��<���<��<r��<L��<Ȝ�<L��<r��<��<���<��<��<���<ا�<���<���<8��<`   `   ���<Ȫ�<���<W��<\��<e��<���<���<��<g��<Ԝ�<���<B��<���<Ԝ�<g��<��<���<���<e��<\��<W��<���<Ȫ�<`   `   ��<��<��<��<p��<x��<��<���<�<d��<���<��<Y��<��<���<d��<�<���<��<x��<p��<��<��<��<`   `   ب�<���<���<	��<Y��<���<��<��<9��<���<ݛ�<���<���<���<ݛ�<���<9��<��<��<���<Y��<	��<���<���<`   `   ���<���<���<���<:��<ݢ�<��<y��<؝�<ԛ�<��<P��<W��<P��<��<ԛ�<؝�<y��<��<ݢ�<:��<���<���<���<`   `   i��<��<}��<���<��<���<���<<��<���<���<u��<���<���<���<u��<���<���<<��<���<���<��<���<}��<��<`   `   E��<���<j��<e��<���<Р�<��<b��<���<���<���<$��<"��<$��<���<���<���<b��<��<Р�<���<e��<j��<���<`   `   ���<`��<(��<��<Ơ�<��<@��<��<ޛ�<���<���<)��<���<)��<���<���<ޛ�<��<@��<��<Ơ�<��<(��<`��<`   `   "��<%��<��<��<��<̞�<e��<���<��<���<���<��<L��<��<���<���<��<���<e��<̞�<��<��<��<%��<`   `   ���<k��<���<P��<^��<o��<j��<���<o��<���<$��<}��<\��<}��<$��<���<o��<���<j��<o��<^��<P��<���<k��<`   `   ���<P��<��<���<��<x��<���<���<��<+��<ך�<j��<H��<j��<ך�<+��<��<���<���<x��<��<���<��<P��<`   `   ��<���<a��<��<���<��<h��<��<���<4��<��<?��<��<?��<��<4��<���<��<h��<��<���<��<a��<���<`   `   ��<F��<��<��<Ȟ�<��<��<ם�<��<���<Ɯ�<���<Ɯ�<���<Ɯ�<���<��<ם�<��<��<Ȟ�<��<��<F��<`   `   Ӟ�<��<Ş�<��<��<���<���<���<��<;��<��<L��<��<L��<��<;��<��<���<���<���<��<��<Ş�<��<`   `   ���<˞�<͞�<���<��<��<l��<\��<���<"��<���<��</��<��<���<"��<���<\��<l��<��<��<���<͞�<˞�<`   `   N��<���<���<.��<f��<̟�<s��<���<��<Y��<���<���<��<���<���<Y��<��<���<s��<̟�<f��<.��<���<���<`   `   ���<��<���<G��<ӟ�<���<X��<ء�<V��<���<\��<ƣ�<ˣ�<ƣ�<\��<���<V��<ء�<X��<���<ӟ�<G��<���<��<`   `   ؞�<��<��<���<���<~��<9��<4��<<��<���<��<\��<H��<\��<��<���<<��<4��<9��<~��<���<���<��<��<`   `   ���<���<_��<��<��<���<ʢ�<��< ��<��<̦�<F��<G��<F��<̦�<��< ��<��<ʢ�<���<��<��<_��<���<`   `   ���<��<p��<0��<f��<N��<���<��<���<��<	��<���<���<���<	��<��<���<��<���<N��<f��<0��<p��<��<`   `   -��<���<d��<T��<���<Т�<a��<��<��<]��<;��<ѩ�<���<ѩ�<;��<]��<��<��<a��<Т�<���<T��<d��<���<`   `   ���<���<7��<^��<���<&��<���<��<���<��<��<���<C��<���<��<��<���<��<���<&��<���<^��<7��<���<`   `   ��<m��<��<���<P��<.��<���<W��<��<z��<8��<���<Z��<���<8��<z��<��<W��<���<.��<P��<���<��<m��<`   `   ���<9��<g��<t��<���<���<���<U��<��<���<ժ�<��<l��<��<ժ�<���<��<U��<���<���<���<t��<g��<9��<`   `   Ȝ�<L��<r��<��<���<��<��<���<ا�<���<���<8��<��<8��<���<���<ا�<���<��<��<���<��<r��<L��<`   `   B��<���<Ԝ�<g��<��<���<���<e��<\��<W��<���<Ȫ�<���<Ȫ�<���<W��<\��<e��<���<���<��<g��<Ԝ�<���<`   `   Y��<��<���<d��<�<���<��<x��<p��<��<��<��<��<��<��<��<p��<x��<��<���<�<d��<���<��<`   `   ���<���<ݛ�<���<9��<��<��<���<Y��<	��<���<���<ب�<���<���<	��<Y��<���<��<��<9��<���<ݛ�<���<`   `   W��<P��<��<ԛ�<؝�<y��<��<ݢ�<:��<���<���<���<���<���<���<���<:��<ݢ�<��<y��<؝�<ԛ�<��<P��<`   `   ���<���<u��<���<���<<��<���<���<��<���<}��<��<i��<��<}��<���<��<���<���<<��<���<���<u��<���<`   `   "��<$��<���<���<���<b��<��<Р�<���<e��<j��<���<E��<���<j��<e��<���<Р�<��<b��<���<���<���<$��<`   `   ���<��<���<���<��<��<��<��<5��<���<-��<Š�<��<Š�<-��<���<5��<��<��<��<��<���<���<��<`   `   ���<���<���<��<���<���<���<|��<O��<���<j��<��<���<��<j��<���<O��<|��<���<���<���<��<���<���<`   `   ؙ�<���<��<T��<њ�<i��<M��<
��<���<K��<���<7��<E��<7��<���<K��<���<
��<M��<i��<њ�<T��<��<���<`   `   ���<��</��<���<C��<���<A��<��<k��<��<��<5��<a��<5��<��<��<k��<��<A��<���<C��<���</��<��<`   `   ֚�<���<��<.��<t��<ʛ�<(��<���<0��<���<Н�<	��<1��<	��<Н�<���<0��<���<(��<ʛ�<t��<.��<��<���<`   `   ƛ�<ě�<���<��<��<~��<���<���<���<)��<h��<ԝ�<�<ԝ�<h��<)��<���<���<���<~��<��<��<���<ě�<`   `   ���<��<��<&��<<��<��<\��<A��<0��<��<@��<i��<���<i��<@��<��<0��<A��<\��<��<<��<&��<��<��<`   `   ���<��<��<��<��<���<���<͝�<���<A��<���<���<1��<���<���<A��<���<͝�<���<���<��<��<��<��<`   `   8��<{��<|��<(��<��<Ş�<M��<5��<֝�<���<u��<>��<d��<>��<u��<���<֝�<5��<M��<Ş�<��<(��<|��<{��<`   `   ��<Ԡ�<���<p��<0��<���<��<���<��<	��<U��<��<f��<��<U��<	��<��<���<��<���<0��<p��<���<Ԡ�<`   `   O��<���<��<v��<ڠ�<*��<���<'��<]��<H��<ʝ�<q��<���<q��<ʝ�<H��<]��<'��<���<*��<ڠ�<v��<��<���<`   `   ���<e��<.��<���<��<5��<���<���<ڞ�<3��<˝�<���<J��<���<˝�<3��<ڞ�<���<���<5��<��<���<.��<e��<`   `   ���<V��<��<���<��<��<��< ��<C��<K��<���<\��<��<\��<���<K��<C��< ��<��<��<��<���<��<V��<`   `   ���<%��<Ѥ�<h��<O��<l��<q��<.��<=��<}��<��<j��<��<j��<��<}��<=��<.��<q��<l��<O��<h��<Ѥ�<%��<`   `   =��<��<���<��<ţ�<���<���<@��<*��<N��<ѝ�<M��<�<M��<ѝ�<N��<*��<@��<���<���<ţ�<��<���<��<`   `   ���<U��<��<"��<'��<���<r��<f��<t��<��<h��<��<c��<��<h��<��<t��<f��<r��<���<'��<"��<��<U��<`   `   ��<���<��<Ѥ�<��<ݢ�<]��<Y��<7��<��<$��<���<��<���<$��<��<7��<Y��<]��<ݢ�<��<Ѥ�<��<���<`   `   ���<M��<��<ݤ�<��<���<*��<��<n��<���<���<��<���<��<���<���<n��<��<*��<���<��<ݤ�<��<M��<`   `   0��<���<���<���<|��<��<͠�<v��<��<>��<��<h��<���<h��<��<>��<��<v��<͠�<��<|��<���<���<���<`   `   ���<.��<���<���<���<���<'��<՞�<y��<v��<���<���<ݚ�<���<���<v��<y��<՞�<'��<���<���<���<���<.��<`   `   ��<���<���<4��<��<��<-��<��<���<���<��<p��<:��<p��<��<���<���<��<-��<��<��<4��<���<���<`   `   ���<ޣ�<b��<f��<j��<@��<���<g��<|��<��<8��<͙�<ҙ�<͙�<8��<��<|��<g��<���<@��<j��<f��<b��<ޣ�<`   `   ���<���<2��<o��<���<s��<*��<��<���<ʚ�<;��<o��<6��<o��<;��<ʚ�<���<��<*��<s��<���<o��<2��<���<`   `   ;��<ǡ�<��<���<���<���<j��<X��<��<^��<$��<=��<̘�<=��<$��<^��<��<X��<j��<���<���<���<��<ǡ�<`   `   ��<Š�<-��<���<5��<��<��<��<��<���<���<��<���<��<���<���<��<��<��<��<5��<���<-��<Š�<`   `   ���<��<j��<���<O��<|��<���<���<���<��<���<���<���<���<���<��<���<���<���<|��<O��<���<j��<��<`   `   E��<7��<���<K��<���<
��<M��<i��<њ�<T��<��<���<ؙ�<���<��<T��<њ�<i��<M��<
��<���<K��<���<7��<`   `   a��<5��<��<��<k��<��<A��<���<C��<���</��<��<���<��</��<���<C��<���<A��<��<k��<��<��<5��<`   `   1��<	��<Н�<���<0��<���<(��<ʛ�<t��<.��<��<���<֚�<���<��<.��<t��<ʛ�<(��<���<0��<���<Н�<	��<`   `   �<ԝ�<h��<)��<���<���<���<~��<��<��<���<ě�<ƛ�<ě�<���<��<��<~��<���<���<���<)��<h��<ԝ�<`   `   ���<i��<@��<��<0��<A��<\��<��<<��<&��<��<��<���<��<��<&��<<��<��<\��<A��<0��<��<@��<i��<`   `   1��<���<���<A��<���<͝�<���<���<��<��<��<��<���<��<��<��<��<���<���<͝�<���<A��<���<���<`   `   d��<>��<u��<���<֝�<5��<M��<Ş�<��<(��<|��<{��<8��<{��<|��<(��<��<Ş�<M��<5��<֝�<���<u��<>��<`   `   f��<��<U��<	��<��<���<��<���<0��<p��<���<Ԡ�<��<Ԡ�<���<p��<0��<���<��<���<��<	��<U��<��<`   `   ���<q��<ʝ�<H��<]��<'��<���<*��<ڠ�<v��<��<���<O��<���<��<v��<ڠ�<*��<���<'��<]��<H��<ʝ�<q��<`   `   J��<���<˝�<3��<ڞ�<���<���<5��<��<���<.��<e��<���<e��<.��<���<��<5��<���<���<ڞ�<3��<˝�<���<`   `   ��<\��<���<K��<C��< ��<��<��<��<���<��<V��<���<V��<��<���<��<��<��< ��<C��<K��<���<\��<`   `   ��<j��<��<}��<=��<.��<q��<l��<O��<h��<Ѥ�<%��<���<%��<Ѥ�<h��<O��<l��<q��<.��<=��<}��<��<j��<`   `   �<M��<ѝ�<N��<*��<@��<���<���<ţ�<��<���<��<=��<��<���<��<ţ�<���<���<@��<*��<N��<ѝ�<M��<`   `   c��<��<h��<��<t��<f��<r��<���<'��<"��<��<U��<���<U��<��<"��<'��<���<r��<f��<t��<��<h��<��<`   `   ��<���<$��<��<7��<Y��<]��<ݢ�<��<Ѥ�<��<���<��<���<��<Ѥ�<��<ݢ�<]��<Y��<7��<��<$��<���<`   `   ���<��<���<���<n��<��<*��<���<��<ݤ�<��<M��<���<M��<��<ݤ�<��<���<*��<��<n��<���<���<��<`   `   ���<h��<��<>��<��<v��<͠�<��<|��<���<���<���<0��<���<���<���<|��<��<͠�<v��<��<>��<��<h��<`   `   ݚ�<���<���<v��<y��<՞�<'��<���<���<���<���<.��<���<.��<���<���<���<���<'��<՞�<y��<v��<���<���<`   `   :��<p��<��<���<���<��<-��<��<��<4��<���<���<��<���<���<4��<��<��<-��<��<���<���<��<p��<`   `   ҙ�<͙�<8��<��<|��<g��<���<@��<j��<f��<b��<ޣ�<���<ޣ�<b��<f��<j��<@��<���<g��<|��<��<8��<͙�<`   `   6��<o��<;��<ʚ�<���<��<*��<s��<���<o��<2��<���<���<���<2��<o��<���<s��<*��<��<���<ʚ�<;��<o��<`   `   ̘�<=��<$��<^��<��<X��<j��<���<���<���<��<ǡ�<;��<ǡ�<��<���<���<���<j��<X��<��<^��<$��<=��<`   `   ���<И�<���<9��<��<t��<V��<��<���<Z��<��<g��<��<g��<��<Z��<���<��<V��<t��<��<9��<���<И�<`   `   ���<���<��<:��<��<k��<h��<ٛ�<���<���<[��<ʝ�<���<ʝ�<[��<���<���<ٛ�<h��<k��<��<:��<��<���<`   `   h��<ǘ�<��<H��<��<S��<��<`��< ��<���<ʜ�<��<�<��<ʜ�<���< ��<`��<��<S��<��<H��<��<ǘ�<`   `   Ř�<���<o��<���<��<���<���<��<���<��<m��<���<t��<���<m��<��<���<��<���<���<��<���<o��<���<`   `    ��<���<��<���<q��<ݚ�<!��<���<}��<���<��<<��<7��<<��<��<���<}��<���<!��<ݚ�<q��<���<��<���<`   `   W��<���<���<���<���<��<%��<���<���<��<ϛ�<���<��<���<ϛ�<��<���<���<%��<��<���<���<���<���<`   `   њ�<f��<u��<\��<���<c��<\��<���<���<��<���<���<ٛ�<���<���<��<���<���<\��<c��<���<\��<u��<f��<`   `   m��<���<^��<ܛ�< ��<3��<��<���<���<ě�<���<f��<՛�<f��<���<ě�<���<���<��<3��< ��<ܛ�<^��<���<`   `   ���<X��<-��<��<���<���<l��<B��<��<���<���<���<��<���<���<���<��<B��<l��<���<���<��<-��<X��<`   `   ���<��<5��<9��<���<l��<��<̜�<u��<��<��<���<ɛ�<���<��<��<u��<̜�<��<l��<���<9��<5��<��<`   `   ���<L��<-��<��<@��<���<���<��<���<@��<��<���<_��<���<��<@��<���<��<���<���<@��<��<-��<L��<`   `   ?��<5��<��<���<@��<���<7��<E��<���<`��<��<Ǜ�<���<Ǜ�<��<`��<���<E��<7��<���<@��<���<��<5��<`   `   &��<-��<��<M��<��<��<?��<���<��<���<
��< ��<��< ��<
��<���<��<���<?��<��<��<M��<��<-��<`   `   ѡ�<Ρ�<\��<���<3��<3��<���<*��<6��<���<��<���<���<���<��<���<6��<*��<���<3��<3��<���<\��<Ρ�<`   `   ��<#��<̡�<���<���<���<��<��<%��<���<ś�<���<՛�<���<ś�<���<%��<��<��<���<���<���<̡�<#��<`   `   L��<���<C��<b��<Ǡ�<���<О�<���<��<���<���<Q��<���<Q��<���<���<��<���<О�<���<Ǡ�<b��<C��<���<`   `   ���<���<��<���<Ϡ�<՟�<��<��<��<��<a��<��<$��<��<a��<��<��<��<��<՟�<Ϡ�<���<��<���<`   `   ���</��<͡�<���<���<���<���<ŝ�<X��<���<d��<͚�<��<͚�<d��<���<X��<ŝ�<���<���<���<���<͡�</��<`   `   ���<��<ޡ�<6��<��<[��<��<'��<��<F��<��<Q��<s��<Q��<��<F��<��<'��<��<[��<��<6��<ޡ�<��<`   `   ܡ�<���<���<���<ʟ�<:��<ǝ�<��<��<���<<��<ř�<ʙ�<ř�<<��<���<��<��<ǝ�<:��<ʟ�<���<���<���<`   `   ��<���<֠�<'��<W��<u��<���<w��<f��<���<
��<���<f��<���<
��<���<f��<w��<���<u��<W��<'��<֠�<���<`   `   {��<}��<
��<y��<���<l��<��<���<w��<b��<���<4��<��<4��<���<b��<w��<���<��<l��<���<y��<
��<}��<`   `   Ɵ�<��<]��<Ȟ�<;��<��<���<f��<u��<��<֘�<ט�<��<ט�<֘�<��<u��<f��<���<��<;��<Ȟ�<]��<��<`   `   Ş�<��<���<��<���<s��<��<���<j��<���<���<���<��<���<���<���<j��<���<��<s��<���<��<���<��<`   `   ��<g��<��<Z��<���<��<V��<t��<��<9��<���<И�<���<И�<���<9��<��<t��<V��<��<���<Z��<��<g��<`   `   ���<ʝ�<[��<���<���<ٛ�<h��<k��<��<:��<��<���<���<���<��<:��<��<k��<h��<ٛ�<���<���<[��<ʝ�<`   `   �<��<ʜ�<���< ��<`��<��<S��<��<H��<��<ǘ�<h��<ǘ�<��<H��<��<S��<��<`��< ��<���<ʜ�<��<`   `   t��<���<m��<��<���<��<���<���<��<���<o��<���<Ř�<���<o��<���<��<���<���<��<���<��<m��<���<`   `   7��<<��<��<���<}��<���<!��<ݚ�<q��<���<��<���< ��<���<��<���<q��<ݚ�<!��<���<}��<���<��<<��<`   `   ��<���<ϛ�<��<���<���<%��<��<���<���<���<���<W��<���<���<���<���<��<%��<���<���<��<ϛ�<���<`   `   ٛ�<���<���<��<���<���<\��<c��<���<\��<u��<f��<њ�<f��<u��<\��<���<c��<\��<���<���<��<���<���<`   `   ՛�<f��<���<ě�<���<���<��<3��< ��<ܛ�<^��<���<m��<���<^��<ܛ�< ��<3��<��<���<���<ě�<���<f��<`   `   ��<���<���<���<��<B��<l��<���<���<��<-��<X��<���<X��<-��<��<���<���<l��<B��<��<���<���<���<`   `   ɛ�<���<��<��<u��<̜�<��<l��<���<9��<5��<��<���<��<5��<9��<���<l��<��<̜�<u��<��<��<���<`   `   _��<���<��<@��<���<��<���<���<@��<��<-��<L��<���<L��<-��<��<@��<���<���<��<���<@��<��<���<`   `   ���<Ǜ�<��<`��<���<E��<7��<���<@��<���<��<5��<?��<5��<��<���<@��<���<7��<E��<���<`��<��<Ǜ�<`   `   ��< ��<
��<���<��<���<?��<��<��<M��<��<-��<&��<-��<��<M��<��<��<?��<���<��<���<
��< ��<`   `   ���<���<��<���<6��<*��<���<3��<3��<���<\��<Ρ�<ѡ�<Ρ�<\��<���<3��<3��<���<*��<6��<���<��<���<`   `   ՛�<���<ś�<���<%��<��<��<���<���<���<̡�<#��<��<#��<̡�<���<���<���<��<��<%��<���<ś�<���<`   `   ���<Q��<���<���<��<���<О�<���<Ǡ�<b��<C��<���<L��<���<C��<b��<Ǡ�<���<О�<���<��<���<���<Q��<`   `   $��<��<a��<��<��<��<��<՟�<Ϡ�<���<��<���<���<���<��<���<Ϡ�<՟�<��<��<��<��<a��<��<`   `   ��<͚�<d��<���<X��<ŝ�<���<���<���<���<͡�</��<���</��<͡�<���<���<���<���<ŝ�<X��<���<d��<͚�<`   `   s��<Q��<��<F��<��<'��<��<[��<��<6��<ޡ�<��<���<��<ޡ�<6��<��<[��<��<'��<��<F��<��<Q��<`   `   ʙ�<ř�<<��<���<��<��<ǝ�<:��<ʟ�<���<���<���<ܡ�<���<���<���<ʟ�<:��<ǝ�<��<��<���<<��<ř�<`   `   f��<���<
��<���<f��<w��<���<u��<W��<'��<֠�<���<��<���<֠�<'��<W��<u��<���<w��<f��<���<
��<���<`   `   ��<4��<���<b��<w��<���<��<l��<���<y��<
��<}��<{��<}��<
��<y��<���<l��<��<���<w��<b��<���<4��<`   `   ��<ט�<֘�<��<u��<f��<���<��<;��<Ȟ�<]��<��<Ɵ�<��<]��<Ȟ�<;��<��<���<f��<u��<��<֘�<ט�<`   `   ��<���<���<���<j��<���<��<s��<���<��<���<��<Ş�<��<���<��<���<s��<��<���<j��<���<���<���<`   `   ��<���<��<���<���<��<͙�<���<ښ�<M��<ɛ�<֛�<��<֛�<ɛ�<M��<ښ�<���<͙�<��<���<���<��<���<`   `   ���<���<���<U��<֘�<��<���<���<m��<��<&��<[��<���<[��<&��<��<m��<���<���<��<֘�<U��<���<���<`   `   ��<��<��<]��<���<��<~��<��<u��<���<���<��<#��<��<���<���<u��<��<~��<��<���<]��<��<��<`   `   ,��<]��<���<Ƙ�<���<��<t��<�<N��<\��<���<Κ�<��<Κ�<���<\��<N��<�<t��<��<���<Ƙ�<���<]��<`   `   ���<���<Ø�<��<��<V��<���<���<��<��<A��<8��<2��<8��<A��<��<��<���<���<V��<��<��<Ø�<���<`   `   a��<��<���<J��<Z��<n��<���<���<���<ޙ�<��<��<"��<��<��<ޙ�<���<���<���<n��<Z��<J��<���<��<`   `   ��<���<���<ݙ�<���<��<��<���<Ù�<ޙ�<$��<U��<���<U��<$��<ޙ�<Ù�<���<��<��<���<ݙ�<���<���<`   `   Ț�<h��<o��<К�<e��<s��<���<B��<1��<$��<��<��<��<��<��<$��<1��<B��<���<s��<e��<К�<o��<h��<`   `   ;��<���<��<l��<՚�<���<���<b��<Y��<3��<Y��<��<���<��<Y��<3��<Y��<b��<���<���<՚�<l��<��<���<`   `   ś�<��<ϛ�<���<c��<:��<���<���<v��<���<c��<S��<ٙ�<S��<c��<���<v��<���<���<:��<c��<���<ϛ�<��<`   `   ���<��<���<A��<=��<ٛ�<K��<���<ߚ�<+��<��<:��<��<:��<��<+��<ߚ�<���<K��<ٛ�<=��<A��<���<��<`   `   (��<D��<��<ל�<���<��<���<D��<%��<���<#��<!��<	��<!��<#��<���<%��<D��<���<��<���<ל�<��<D��<`   `   ܝ�<ܝ�<���<P��<��<~��<��<���<���<���<P��<��<��<��<P��<���<���<���<��<~��<��<P��<���<ܝ�<`   `   ���<p��<^��<���<���<���<*��<���<��<���<B��<��<ș�<��<B��<���<��<���<*��<���<���<���<^��<p��<`   `   ��<Ξ�<a��<G��<Ν�<��<M��<ߛ�<��<���<\��<ߙ�<���<ߙ�<\��<���<��<ߛ�<M��<��<Ν�<G��<a��<Ξ�<`   `   <��<��<|��<`��<���<ʜ�<���<Û�<��<���<k��<ə�<���<ə�<k��<���<��<Û�<���<ʜ�<���<`��<|��<��<`   `   ̞�<'��<���<���<���<��<o��<g��<ך�<F��<���<~��<���<~��<���<F��<ך�<g��<o��<��<���<���<���<'��<`   `   ��<H��<���<A��<x��<���<5��<k��<��<��<���<5��<A��<5��<���<��<��<k��<5��<���<x��<A��<���<H��<`   `   ���<��<]��<���<E��<ڜ�<ڛ�< ��<���<˙�<~��<��<ј�<��<~��<˙�<���< ��<ڛ�<ڜ�<E��<���<]��<��<`   `   5��<}��<*��<~��<��<P��<^��<���<���<T��<��<���<���<���<��<T��<���<���<^��<P��<��<~��<*��<}��<`   `   L��<&��<���<6��<Ŝ�<˛�<C��<���<���<��<���<���<Z��<���<���<��<���<���<C��<˛�<Ŝ�<6��<���<&��<`   `   ��<o��<��<���<V��<b��<��<S��<���<��<x��<O��<���<O��<x��<��<���<S��<��<b��<V��<���<��<o��<`   `   ^��<��<���<C��<ޛ�<!��<@��<���<-��<���<3��<��<���<��<3��<���<-��<���<@��<!��<ޛ�<C��<���<��<`   `   ���<U��<b��<���<|��<��<��<`��<͘�<i��<��<ϗ�<V��<ϗ�<��<i��<͘�<`��<��<��<|��<���<b��<U��<`   `   ��<֛�<ɛ�<M��<ښ�<���<͙�<��<���<���<��<���<��<���<��<���<���<��<͙�<���<ښ�<M��<ɛ�<֛�<`   `   ���<[��<&��<��<m��<���<���<��<֘�<U��<���<���<���<���<���<U��<֘�<��<���<���<m��<��<&��<[��<`   `   #��<��<���<���<u��<��<~��<��<���<]��<��<��<��<��<��<]��<���<��<~��<��<u��<���<���<��<`   `   ��<Κ�<���<\��<N��<�<t��<��<���<Ƙ�<���<]��<,��<]��<���<Ƙ�<���<��<t��<�<N��<\��<���<Κ�<`   `   2��<8��<A��<��<��<���<���<V��<��<��<Ø�<���<���<���<Ø�<��<��<V��<���<���<��<��<A��<8��<`   `   "��<��<��<ޙ�<���<���<���<n��<Z��<J��<���<��<a��<��<���<J��<Z��<n��<���<���<���<ޙ�<��<��<`   `   ���<U��<$��<ޙ�<Ù�<���<��<��<���<ݙ�<���<���<��<���<���<ݙ�<���<��<��<���<Ù�<ޙ�<$��<U��<`   `   ��<��<��<$��<1��<B��<���<s��<e��<К�<o��<h��<Ț�<h��<o��<К�<e��<s��<���<B��<1��<$��<��<��<`   `   ���<��<Y��<3��<Y��<b��<���<���<՚�<l��<��<���<;��<���<��<l��<՚�<���<���<b��<Y��<3��<Y��<��<`   `   ٙ�<S��<c��<���<v��<���<���<:��<c��<���<ϛ�<��<ś�<��<ϛ�<���<c��<:��<���<���<v��<���<c��<S��<`   `   ��<:��<��<+��<ߚ�<���<K��<ٛ�<=��<A��<���<��<���<��<���<A��<=��<ٛ�<K��<���<ߚ�<+��<��<:��<`   `   	��<!��<#��<���<%��<D��<���<��<���<ל�<��<D��<(��<D��<��<ל�<���<��<���<D��<%��<���<#��<!��<`   `   ��<��<P��<���<���<���<��<~��<��<P��<���<ܝ�<ܝ�<ܝ�<���<P��<��<~��<��<���<���<���<P��<��<`   `   ș�<��<B��<���<��<���<*��<���<���<���<^��<p��<���<p��<^��<���<���<���<*��<���<��<���<B��<��<`   `   ���<ߙ�<\��<���<��<ߛ�<M��<��<Ν�<G��<a��<Ξ�<��<Ξ�<a��<G��<Ν�<��<M��<ߛ�<��<���<\��<ߙ�<`   `   ���<ə�<k��<���<��<Û�<���<ʜ�<���<`��<|��<��<<��<��<|��<`��<���<ʜ�<���<Û�<��<���<k��<ə�<`   `   ���<~��<���<F��<ך�<g��<o��<��<���<���<���<'��<̞�<'��<���<���<���<��<o��<g��<ך�<F��<���<~��<`   `   A��<5��<���<��<��<k��<5��<���<x��<A��<���<H��<��<H��<���<A��<x��<���<5��<k��<��<��<���<5��<`   `   ј�<��<~��<˙�<���< ��<ڛ�<ڜ�<E��<���<]��<��<���<��<]��<���<E��<ڜ�<ڛ�< ��<���<˙�<~��<��<`   `   ���<���<��<T��<���<���<^��<P��<��<~��<*��<}��<5��<}��<*��<~��<��<P��<^��<���<���<T��<��<���<`   `   Z��<���<���<��<���<���<C��<˛�<Ŝ�<6��<���<&��<L��<&��<���<6��<Ŝ�<˛�<C��<���<���<��<���<���<`   `   ���<O��<x��<��<���<S��<��<b��<V��<���<��<o��<��<o��<��<���<V��<b��<��<S��<���<��<x��<O��<`   `   ���<��<3��<���<-��<���<@��<!��<ޛ�<C��<���<��<^��<��<���<C��<ޛ�<!��<@��<���<-��<���<3��<��<`   `   V��<ϗ�<��<i��<͘�<`��<��<��<|��<���<b��<U��<���<U��<b��<���<|��<��<��<`��<͘�<i��<��<ϗ�<`   `   ��<���<��<��<��<!��<2��<���<*��<��<~��<���<��<���<~��<��<*��<���<2��<!��<��<��<��<���<`   `   ���<���<���<��<��<���<̗�<M��<���<��<n��<J��<���<J��<n��<��<���<M��<̗�<���<��<��<���<���<`   `   ɖ�<̖�<ʖ�<��<L��<���<���<Q��<8��<���<��<��<���<��<��<���<8��<Q��<���<���<L��<��<ʖ�<̖�<`   `   ���<��<Ֆ�<(��<I��<���<��<��<:��<m��<���<���<ј�<���<���<m��<:��<��<��<���<I��<(��<Ֆ�<��<`   `   ��<��<��<g��<���<ɗ�<��<��<g��<���<���<���<Ә�<���<���<���<g��<��<��<ɗ�<���<g��<��<��<`   `   ���<ؗ�<��<��<��<��<��<.��<t��<c��<}��<~��<c��<~��<}��<c��<t��<.��<��<��<��<��<��<ؗ�<`   `   (��<?��<t��<��<��<E��<'��<b��<s��<��<<��<>��<ԗ�<>��<<��<��<s��<b��<'��<E��<��<��<t��<?��<`   `   u��<r��<���<{��<���<h��<9��<b��<���<7��<.��<b��<7��<b��<.��<7��<���<b��<9��<h��<���<{��<���<r��<`   `   3��<m��<*��<��<#��<���<���<���<���<���<,��<b��<���<b��<,��<���<���<���<���<���<#��<��<*��<m��<`   `   ���<!��<���<A��<|��<Q��<W��<͘�<���<���<��<���<C��<���<��<���<���<͘�<W��<Q��<|��<A��<���<!��<`   `   ��<i��<'��<��<��<���<O��<��<ј�<ʘ�<y��<D��<c��<D��<y��<ʘ�<ј�<��<O��<���<��<��<'��<i��<`   `    ��<ݚ�<���<̚�<5��<���<���<A��<ݘ�<���<���<a��<O��<a��<���<���<ݘ�<A��<���<���<5��<̚�<���<ݚ�<`   `   ���<C��<��<ߚ�<W��<^��<��<���<���<���<���<E��<#��<E��<���<���<���<���<��<^��<W��<ߚ�<��<C��<`   `   ���<X��<w��<��<���<���<��<Q��<B��<ژ�<���<���<}��<���<���<ژ�<B��<Q��<��<���<���<��<w��<X��<`   `   ��<���<�<u��<���<r��<ș�<r��<W��<���<Z��<b��<8��<b��<Z��<���<W��<r��<ș�<r��<���<u��<�<���<`   `   3��<��<���<���<'��<̚�<B��<ř�<2��<Y��<E��<��<ח�<��<E��<Y��<2��<ř�<B��<̚�<'��<���<���<��<`   `   ��<+��<���<j��<B��<ښ�<���<X��<)��<~��<T��<��<���<��<T��<~��<)��<X��<���<ښ�<B��<j��<���<+��<`   `   ���<F��<���<n��<���<_��<���<���<��<>��<���<ۗ�<ї�<ۗ�<���<>��<��<���<���<_��<���<n��<���<F��<`   `   ���<ӛ�<k��<���<��<:��<-��<;��<���<��<ח�<���<o��<���<ח�<��<���<;��<-��<:��<��<���<k��<ӛ�<`   `   ���<���<4��<O��<���<���<���<��<J��<E��<���<M��<D��<M��<���<E��<J��<��<���<���<���<O��<4��<���<`   `   ���<a��<&��<���<D��<���<"��<~��<7��<��<��<���<��<���<��<��<7��<~��<"��<���<D��<���<&��<a��<`   `   ���<���<��<o��<��<���<��<X��<��<n��<��<���<ږ�<���<��<n��<��<X��<��<���<��<o��<��<���<`   `   ���<S��<���<��<C��<,��<R��<��<���<!��<��<ߖ�<���<ߖ�<��<!��<���<��<R��<,��<C��<��<���<S��<`   `   ���<���<��<���<��<���<W��<Q��<c��<��<��<���<Ֆ�<���<��<��<c��<Q��<W��<���<��<���<��<���<`   `   ��<���<~��<��<*��<���<2��<!��<��<��<��<���<��<���<��<��<��<!��<2��<���<*��<��<~��<���<`   `   ���<J��<n��<��<���<M��<̗�<���<��<��<���<���<���<���<���<��<��<���<̗�<M��<���<��<n��<J��<`   `   ���<��<��<���<8��<Q��<���<���<L��<��<ʖ�<̖�<ɖ�<̖�<ʖ�<��<L��<���<���<Q��<8��<���<��<��<`   `   ј�<���<���<m��<:��<��<��<���<I��<(��<Ֆ�<��<���<��<Ֆ�<(��<I��<���<��<��<:��<m��<���<���<`   `   Ә�<���<���<���<g��<��<��<ɗ�<���<g��<��<��<��<��<��<g��<���<ɗ�<��<��<g��<���<���<���<`   `   c��<~��<}��<c��<t��<.��<��<��<��<��<��<ؗ�<���<ؗ�<��<��<��<��<��<.��<t��<c��<}��<~��<`   `   ԗ�<>��<<��<��<s��<b��<'��<E��<��<��<t��<?��<(��<?��<t��<��<��<E��<'��<b��<s��<��<<��<>��<`   `   7��<b��<.��<7��<���<b��<9��<h��<���<{��<���<r��<u��<r��<���<{��<���<h��<9��<b��<���<7��<.��<b��<`   `   ���<b��<,��<���<���<���<���<���<#��<��<*��<m��<3��<m��<*��<��<#��<���<���<���<���<���<,��<b��<`   `   C��<���<��<���<���<͘�<W��<Q��<|��<A��<���<!��<���<!��<���<A��<|��<Q��<W��<͘�<���<���<��<���<`   `   c��<D��<y��<ʘ�<ј�<��<O��<���<��<��<'��<i��<��<i��<'��<��<��<���<O��<��<ј�<ʘ�<y��<D��<`   `   O��<a��<���<���<ݘ�<A��<���<���<5��<̚�<���<ݚ�< ��<ݚ�<���<̚�<5��<���<���<A��<ݘ�<���<���<a��<`   `   #��<E��<���<���<���<���<��<^��<W��<ߚ�<��<C��<���<C��<��<ߚ�<W��<^��<��<���<���<���<���<E��<`   `   }��<���<���<ژ�<B��<Q��<��<���<���<��<w��<X��<���<X��<w��<��<���<���<��<Q��<B��<ژ�<���<���<`   `   8��<b��<Z��<���<W��<r��<ș�<r��<���<u��<�<���<��<���<�<u��<���<r��<ș�<r��<W��<���<Z��<b��<`   `   ח�<��<E��<Y��<2��<ř�<B��<͚�<'��<���<���<��<3��<��<���<���<'��<͚�<B��<ř�<2��<Y��<E��<��<`   `   ���<��<T��<~��<)��<X��<���<ښ�<B��<j��<���<+��<��<+��<���<j��<B��<ښ�<���<X��<)��<~��<T��<��<`   `   ї�<ۗ�<���<>��<��<���<���<_��<���<n��<���<F��<���<F��<���<n��<���<_��<���<���<��<>��<���<ۗ�<`   `   o��<���<ח�<��<���<;��<-��<:��<��<���<k��<ӛ�<���<ӛ�<k��<���<��<:��<-��<;��<���<��<ח�<���<`   `   D��<M��<���<E��<J��<��<���<���<���<O��<4��<���<���<���<4��<O��<���<���<���<��<J��<E��<���<M��<`   `   ��<���<��<��<7��<~��<"��<���<D��<���<&��<a��<���<a��<&��<���<D��<���<"��<~��<7��<��<��<���<`   `   ږ�<���<��<n��<��<X��<��<���<��<o��<��<���<���<���<��<o��<��<���<��<X��<��<n��<��<���<`   `   ���<ߖ�<��<!��<���<��<R��<,��<C��<��<���<S��<���<S��<���<��<C��<,��<R��<��<���<!��<��<ߖ�<`   `   Ֆ�<���<��<��<c��<Q��<W��<���<��<���<��<���<���<���<��<���<��<���<W��<Q��<c��<��<��<���<`   `   {��<3��<T��<���<	��<	��<Z��<���<��<.��<y��<ɗ�<E��<ɗ�<y��<.��<��<���<Z��<	��<	��<���<T��<3��<`   `   ��<X��<���<���<��<��<G��<Ȗ�<��<��<;��<o��<K��<o��<;��<��<��<Ȗ�<G��<��<��<���<���<X��<`   `   ��<Y��<���<ƕ�<���<*��<<��<���<��< ��<2��<2��<G��<2��<2��< ��<��<���<<��<*��<���<ƕ�<���<Y��<`   `   ���<ە�<ȕ�<��<��<$��<%��<d��<���<Ė�<���<��<��<��<���<Ė�<���<d��<%��<$��<��<��<ȕ�<ە�<`   `   ���<&��<��<��<��<��<f��<���<i��<n��<���<���<ٖ�<���<���<n��<i��<���<f��<��<��<��<��<&��<`   `   ���<��<��<��<K��<4��<v��<���<j��<���<���<���<��<���<���<���<j��<���<v��<4��<K��<��<��<��<`   `   s��<M��<b��<U��<���<���<h��<n��<���<ݖ�<���<���<y��<���<���<ݖ�<���<n��<h��<���<���<U��<b��<M��<`   `   ��<��<��<���<��<���<Ζ�<���<���<���<���<���<���<���<���<���<���<���<Ζ�<���<��<���<��<��<`   `   X��<_��<T��<��<9��<��<��<���<���<���<���<���<���<���<���<���<���<���<��<��<9��<��<T��<_��<`   `   ���<���<���<���<x��<��<��<��<Ֆ�<ږ�<���<���<���<���<���<ږ�<Ֆ�<��<��<��<x��<���<���<���<`   `   ��<ܗ�<��<���<~��<���<e��<6��<��<ǖ�<ޖ�<���<���<���<ޖ�<ǖ�<��<6��<e��<���<~��<���<��<ܗ�<`   `   d��<J��<J��<,��<��<��<���<[��<���<���<ǖ�<���<���<���<ǖ�<���<���<[��<���<��<��<,��<J��<J��<`   `   ���<���<���<���<u��<ڗ�<R��<i��<1��<��<���<���<���<���<���<��<1��<i��<R��<ڗ�<u��<���<���<���<`   `   ��<)��<��<���<���<��<ԗ�<���<K��<��<���<���<���<���<���<��<K��<���<ԗ�<��<���<���<��<)��<`   `   I��<M��<6��<Ø�<���<c��<"��<}��<��<��<���<���<o��<���<���<��<��<}��<"��<c��<���<Ø�<6��<M��<`   `   V��<N��<f��<��<���<9��<���<^��<���<���<���<���<���<���<���<���<���<^��<���<9��<���<��<f��<N��<`   `   e��<D��<T��<��<���<:��<ח�<���<��<���<���<A��<a��<A��<���<���<��<���<ח�<:��<���<��<T��<D��<`   `   n��<:��<:��<ߘ�<j��<��<ї�<��<ٖ�<���<u��</��<*��</��<u��<���<ٖ�<��<ї�<��<j��<ߘ�<:��<:��<`   `   m��<6��<��<Ƙ�<B��<��<���<%��<���<X��<��<%��<!��<%��<��<X��<���<%��<���<��<B��<Ƙ�<��<6��<`   `   /��<��<��<{��<5��<��<}��<(��<���<F��<���<��<��<��<���<F��<���<(��<}��<��<5��<{��<��<��<`   `   Ř�<�<���</��<��<���</��<��<T��<��<��<͕�<˕�<͕�<��<��<T��<��</��<���<��</��<���<�<`   `   ���<���<S��<��<���<z��<!��<���<��<��<��<���<���<���<��<��<��<���<!��<z��<���<��<S��<���<`   `   ��<j��<���<���<���<A��<	��<g��< ��< ��<���<>��<v��<>��<���< ��< ��<g��<	��<A��<���<���<���<j��<`   `   ���<��<���<���<x��<��<���<"��<��<��<=��<��<V��<��<=��<��<��<"��<���<��<x��<���<���<��<`   `   E��<ɗ�<y��<.��<��<���<Z��<	��<	��<���<T��<3��<{��<3��<T��<���<	��<	��<Z��<���<��<.��<y��<ɗ�<`   `   K��<o��<;��<��<��<Ȗ�<G��<��<��<���<���<X��<��<X��<���<���<��<��<G��<Ȗ�<��<��<;��<o��<`   `   G��<2��<2��< ��<��<���<<��<*��<���<ƕ�<���<Y��<��<Y��<���<ƕ�<���<*��<<��<���<��< ��<2��<2��<`   `   ��<��<���<Ė�<���<d��<%��<$��<��<��<ȕ�<ە�<���<ە�<ȕ�<��<��<$��<%��<d��<���<Ė�<���<��<`   `   ٖ�<���<���<n��<i��<���<f��<��<��<��<��<&��<���<&��<��<��<��<��<f��<���<i��<n��<���<���<`   `   ��<���<���<���<j��<���<v��<4��<K��<��<��<��<���<��<��<��<K��<4��<v��<���<j��<���<���<���<`   `   y��<���<���<ݖ�<���<n��<h��<���<���<U��<b��<M��<s��<M��<b��<U��<���<���<h��<n��<���<ݖ�<���<���<`   `   ���<���<���<���<���<���<Ζ�<���<��<���<��<��<��<��<��<���<��<���<Ζ�<���<���<���<���<���<`   `   ���<���<���<���<���<���<��<��<9��<��<T��<_��<X��<_��<T��<��<9��<��<��<���<���<���<���<���<`   `   ���<���<���<ږ�<Ֆ�<��<��<��<x��<���<���<���<���<���<���<���<x��<��<��<��<Ֆ�<ږ�<���<���<`   `   ���<���<ޖ�<ǖ�<��<6��<e��<���<~��<���<��<ܗ�<��<ܗ�<��<���<~��<���<e��<6��<��<ǖ�<ޖ�<���<`   `   ���<���<ǖ�<���<���<[��<���<��<��<,��<J��<J��<d��<J��<J��<,��<��<��<���<[��<���<���<ǖ�<���<`   `   ���<���<���<��<1��<i��<R��<ڗ�<u��<���<���<���<���<���<���<���<u��<ڗ�<R��<i��<1��<��<���<���<`   `   ���<���<���<��<K��<���<ԗ�<��<���<���<��<)��<��<)��<��<���<���<��<ԗ�<���<K��<��<���<���<`   `   o��<���<���<��<��<}��<"��<c��<���<Ø�<6��<M��<I��<M��<6��<Ø�<���<c��<"��<}��<��<��<���<���<`   `   ���<���<���<���<���<^��<���<9��<���<��<f��<N��<V��<N��<f��<��<���<9��<���<^��<���<���<���<���<`   `   a��<A��<���<���<��<���<ח�<:��<���<��<T��<D��<e��<D��<T��<��<���<:��<ח�<���<��<���<���<A��<`   `   *��</��<u��<���<ٖ�<��<ї�<��<j��<ߘ�<:��<:��<n��<:��<:��<ߘ�<j��<��<ї�<��<ٖ�<���<u��</��<`   `   !��<%��<��<X��<���<%��<���<��<B��<Ƙ�<��<6��<m��<6��<��<Ƙ�<B��<��<���<%��<���<X��<��<%��<`   `   ��<��<���<F��<���<(��<}��<��<5��<{��<��<��</��<��<��<{��<5��<��<}��<(��<���<F��<���<��<`   `   ˕�<͕�<��<��<T��<��</��<���<��</��<���<�<Ř�<�<���</��<��<���</��<��<T��<��<��<͕�<`   `   ���<���<��<��<��<���<!��<z��<���<��<S��<���<���<���<S��<��<���<z��<!��<���<��<��<��<���<`   `   v��<>��<���< ��< ��<g��<	��<A��<���<���<���<j��<��<j��<���<���<���<A��<	��<g��< ��< ��<���<>��<`   `   V��<��<=��<��<��<"��<���<��<x��<���<���<��<���<��<���<���<x��<��<���<"��<��<��<=��<��<`   `   ���<��<��<���<���<i��<��<	��<��<���<���<��<���<��<���<���<��<	��<��<i��<���<���<��<��<`   `   (��<'��<��<���<o��<���<���<��<���<_��<%��<j��<���<j��<%��<_��<���<��<���<���<o��<���<��<'��<`   `   ���<��<Γ�<���<��<w��<���<���<���<,��<��<0��<}��<0��<��<,��<���<���<���<w��<��<���<Γ�<��<`   `   2��<���<��<H��<?��<���<���<���<
��<
��<,��<I��<6��<I��<,��<
��<
��<���<���<���<?��<H��<��<���<`   `   #��<H��<t��<���<���<���<���<��<���<��<4��<��<���<��<4��<��<���<��<���<���<���<���<t��<H��<`   `   ���<z��<r��<���<���<���<ʔ�<Ŕ�<���<��<��<��<���<��<��<��<���<Ŕ�<ʔ�<���<���<���<r��<z��<`   `   1��<���<Δ�<��<��<���<��<��<ɔ�<��<���<���<B��<���<���<��<ɔ�<��<��<���<��<��<Δ�<���<`   `   >��<���<\��<N��<��<۔�<��<!��<��<��<���<ٔ�<���<ٔ�<���<��<��<!��<��<۔�<��<N��<\��<���<`   `   =��<��<W��<+��<��<(��<��<��<
��<��<��<Ĕ�<T��<Ĕ�<��<��<
��<��<��<(��<��<+��<W��<��<`   `   ��<���<���<���<���<s��<���<��<.��<ޔ�<��<��<�<��<��<ޔ�<.��<��<���<s��<���<���<���<���<`   `   ���<3��<��<��<���<ʕ�<M��<E��<D��<Ô�<��<��<���<��<��<Ô�<D��<E��<M��<ʕ�<���<��<��<3��<`   `   8��<h��<P��<Ε�<Õ�<%��<���<p��<y��<2��<���<���<Δ�<���<���<2��<y��<p��<���<%��<Õ�<Ε�<P��<h��<`   `    ��<���<t��<4��<7��<Ǖ�<���<l��<I��<W��<-��<��<��<��<-��<W��<I��<l��<���<Ǖ�<7��<4��<t��<���<`   `   ���<ז�<z��<}��<h��<���< ��<���<���<��<���<���<���<���<���<��<���<���< ��<���<h��<}��<z��<ז�<`   `   ږ�<���<���<���<���<��<'��<���<@��<4��<��<���<z��<���<��<4��<@��<���<'��<��<���<���<���<���<`   `   ��<�<Ȗ�<���<m��<��<���<���<P��<S��<��<���<���<���<��<S��<P��<���<���<��<m��<���<Ȗ�<�<`   `   j��<ږ�<��<���<w��<��<ܕ�<ŕ�<���<��<���<���<���<���<���<��<���<ŕ�<ܕ�<��<w��<���<��<ږ�<`   `   !��<���<��<���<���<b��<ߕ�<���<��<��<ؔ�<���<}��<���<ؔ�<��<��<���<ߕ�<b��<���<���<��<���<`   `   ��<���<Ԗ�<J��<E��<.��<D��<,��<\��<��<���<���<X��<���<���<��<\��<,��<D��<.��<E��<J��<Ԗ�<���<`   `   ���<���<���<G��<G��<2��<X��<1��<��<���<l��<a��<"��<a��<l��<���<��<1��<X��<2��<G��<G��<���<���<`   `   n��<m��<���<~��<=��<ŕ�<G��</��<ɔ�<x��<���<8��<
��<8��<���<x��<ɔ�</��<G��<ŕ�<=��<~��<���<m��<`   `   ���<v��<��<+��<ŕ�<��<��<��<ה�<h��<(��<Փ�<��<Փ�<(��<h��<ה�<��<��<��<ŕ�<+��<��<v��<`   `   Օ�<,��<���<ܕ�<���</��<4��<Ӕ�<���<7��<6��<+��<%��<+��<6��<7��<���<Ӕ�<4��</��<���<ܕ�<���<,��<`   `   b��<��<���<���<���<5��<#��<a��<p��<	��<c��<d��<��<d��<c��<	��<p��<a��<#��<5��<���<���<���<��<`   `   ���<��<���<���<��<	��<��<i��<���<���<��<��<���<��<��<���<���<i��<��<	��<��<���<���<��<`   `   ���<j��<%��<_��<���<��<���<���<o��<���<��<'��<(��<'��<��<���<o��<���<���<��<���<_��<%��<j��<`   `   }��<0��<��<,��<���<���<���<w��<��<���<Γ�<��<���<��<Γ�<���<��<w��<���<���<���<,��<��<0��<`   `   6��<I��<,��<
��<
��<���<���<���<?��<H��<��<���<2��<���<��<H��<?��<���<���<���<
��<
��<,��<I��<`   `   ���<��<4��<��<���<��<���<���<���<���<t��<H��<#��<H��<t��<���<���<���<���<��<���<��<4��<��<`   `   ���<��<��<��<���<Ŕ�<ʔ�<���<���<���<r��<z��<���<z��<r��<���<���<���<ʔ�<Ŕ�<���<��<��<��<`   `   B��<���<���<��<ɔ�<��<��<���<��<��<Δ�<���<1��<���<Δ�<��<��<���<��<��<ɔ�<��<���<���<`   `   ���<ٔ�<���<��<��<!��<��<۔�<��<N��<\��<���<>��<���<\��<N��<��<۔�<��<!��<��<��<���<ٔ�<`   `   T��<Ĕ�<��<��<
��<��<��<(��<��<+��<W��<��<=��<��<W��<+��<��<(��<��<��<
��<��<��<Ĕ�<`   `   �<��<��<ޔ�<.��<��<���<s��<���<���<���<���<��<���<���<���<���<s��<���<��<.��<ޔ�<��<��<`   `   ���<��<��<Ô�<D��<E��<M��<ʕ�<���<��<��<3��<���<3��<��<��<���<ʕ�<M��<E��<D��<Ô�<��<��<`   `   Δ�<���<���<2��<y��<p��<���<%��<Õ�<Ε�<P��<h��<8��<h��<P��<Ε�<Õ�<%��<���<p��<y��<2��<���<���<`   `   ��<��<-��<W��<I��<l��<���<Ǖ�<7��<4��<t��<���< ��<���<t��<4��<7��<Ǖ�<���<l��<I��<W��<-��<��<`   `   ���<���<���<��<���<���< ��<���<h��<}��<z��<ז�<���<ז�<z��<}��<h��<���< ��<���<���<��<���<���<`   `   z��<���<��<4��<@��<���<'��<��<���<���<���<���<ږ�<���<���<���<���<��<'��<���<@��<4��<��<���<`   `   ���<���<��<S��<P��<���<���<��<m��<���<Ȗ�<�<��<�<Ȗ�<���<m��<��<���<���<P��<S��<��<���<`   `   ���<���<���<��<���<ŕ�<ܕ�<��<w��<���<��<ږ�<j��<ږ�<��<���<w��<��<ܕ�<ŕ�<���<��<���<���<`   `   }��<���<ؔ�<��<��<���<ߕ�<b��<���<���<��<���<!��<���<��<���<���<b��<ߕ�<���<��<��<ؔ�<���<`   `   X��<���<���<��<\��<,��<D��<.��<E��<J��<Ԗ�<���<��<���<Ԗ�<J��<E��<.��<D��<,��<\��<��<���<���<`   `   "��<a��<l��<���<��<1��<X��<2��<G��<G��<���<���<���<���<���<G��<G��<2��<X��<1��<��<���<l��<a��<`   `   
��<8��<���<x��<ɔ�</��<G��<ŕ�<=��<~��<���<m��<n��<m��<���<~��<=��<ŕ�<G��</��<ɔ�<x��<���<8��<`   `   ��<Փ�<(��<h��<ה�<��<��<��<ŕ�<+��<��<v��<���<v��<��<+��<ŕ�<��<��<��<ה�<h��<(��<Փ�<`   `   %��<+��<6��<7��<���<Ӕ�<4��</��<���<ܕ�<���<,��<Օ�<,��<���<ܕ�<���</��<4��<Ӕ�<���<7��<6��<+��<`   `   ��<d��<c��<	��<p��<a��<#��<5��<���<���<���<��<b��<��<���<���<���<5��<#��<a��<p��<	��<c��<d��<`   `   O��<V��<���<���<��<��<��<I��<{��<���<t��<���<��<���<t��<���<{��<I��<��<��<��<���<���<V��<`   `   t��<Y��<���<��<ڒ�<ϒ�<��<I��<v��<ɓ�<œ�<���<���<���<œ�<ɓ�<v��<I��<��<ϒ�<ڒ�<��<���<Y��<`   `   ���<z��<��<��<ߒ�<��<��<5��<!��<Z��<���<���<a��<���<���<Z��<!��<5��<��<��<ߒ�<��<��<z��<`   `   ���<���<ʒ�<��<Ւ�<��<*��<@��< ��<���<<��<g��<\��<g��<<��<���< ��<@��<*��<��<Ւ�<��<ʒ�<���<`   `   ���<В�<��<Ӓ�<��<��<���<��<F��<1��<B��<k��<i��<k��<B��<1��<F��<��<���<��<��<Ӓ�<��<В�<`   `   ��<��<"��<֒�<���<B��<��<��<M��<A��<C��<:��<��<:��<C��<A��<M��<��<��<B��<���<֒�<"��<��<`   `   ��<��<��<��<	��<K��<9��<C��<Q��<)��<>��<)��<��<)��<>��<)��<Q��<C��<9��<K��<	��<��<��<��<`   `   ;��<@��<7��<7��<X��<H��<��<��<@��<7��<R��<g��<Q��<g��<R��<7��<@��<��<��<H��<X��<7��<7��<@��<`   `   ���<ړ�<���<T��<���<���<i��<'��<G��<L��<��<P��<{��<P��<��<L��<G��<'��<i��<���<���<T��<���<ړ�<`   `   ���<���<ԓ�<���<���<ԓ�<��<���<f��<f��<��<,��<b��<,��<��<f��<f��<���<��<ԓ�<���<���<ԓ�<���<`   `   ���<���<Г�<���<ӓ�<o��<���<���<T��<i��<I��<5��<>��<5��<I��<i��<T��<���<���<o��<ӓ�<���<Г�<���<`   `   %��<��<	��<I��<
��<���<���<z��<I��<O��<M��<6��<0��<6��<M��<O��<I��<z��<���<���<
��<I��<	��<��<`   `   ���<w��<H��<`��<"��<'��<��<���<���<X��<3��<4��<7��<4��<3��<X��<���<���<��<'��<"��<`��<H��<w��<`   `   ���<���<x��<^��<��<��<ݓ�<���<ē�<d��<,��<K��<?��<K��<,��<d��<ē�<���<ݓ�<��<��<^��<x��<���<`   `   ���<���<ɔ�<���<(��<*��<���<���<ݓ�<J��<��<R��<*��<R��<��<J��<ݓ�<���<���<*��<(��<���<ɔ�<���<`   `   ���<���<Ҕ�<���<k��<���<��<œ�<Γ�<?��<��<0��<��<0��<��<?��<Γ�<œ�<��<���<k��<���<Ҕ�<���<`   `   Ô�<���<���<N��<7��<!��<��<���<|��<I��<&��<>��<���<>��<&��<I��<|��<���<��<!��<7��<N��<���<���<`   `   ���<���<���<k��<>��<ԓ�<�<y��<M��<7��<��<<��<��<<��<��<7��<M��<y��<�<ԓ�<>��<k��<���<���<`   `   ���<���<���<���<5��<���<���<���<7��<��<͒�<��<ג�<��<͒�<��<7��<���<���<���<5��<���<���<���<`   `   Ҕ�<���<Z��<Z��<���<���<��<���<��<���<��<ݒ�<Ԓ�<ݒ�<��<���<��<���<��<���<���<Z��<Z��<���<`   `   ���<b��<,��<��<œ�<͓�<͓�<+��<��<,��<��<ޒ�<��<ޒ�<��<,��<��<+��<͓�<͓�<œ�<��<,��<b��<`   `   &��<R��<T��<��<˓�<��<���<��<��<���<���<���<��<���<���<���<��<��<���<��<˓�<��<T��<R��<`   `   ���<8��<O��<ߓ�<���<�<K��<
��<��<���<��<}��<���<}��<��<���<��<
��<K��<�<���<ߓ�<O��<8��<`   `   -��<��<�<���<d��<F��<"��<0��<���<���<���<x��<M��<x��<���<���<���<0��<"��<F��<d��<���<�<��<`   `   ��<���<t��<���<{��<I��<��<��<��<���<���<V��<O��<V��<���<���<��<��<��<I��<{��<���<t��<���<`   `   ���<���<œ�<ɓ�<v��<I��<��<ϒ�<ڒ�<��<���<Y��<t��<Y��<���<��<ڒ�<ϒ�<��<I��<v��<ɓ�<œ�<���<`   `   a��<���<���<Z��<!��<5��<��<��<ߒ�<��<��<z��<���<z��<��<��<ߒ�<��<��<5��<!��<Z��<���<���<`   `   \��<g��<<��<���< ��<@��<*��<��<Ւ�<��<ʒ�<���<���<���<ʒ�<��<Ւ�<��<*��<@��< ��<���<<��<g��<`   `   i��<k��<B��<1��<F��<��<���<��<��<Ӓ�<��<В�<���<В�<��<Ӓ�<��<��<���<��<F��<1��<B��<k��<`   `   ��<:��<C��<A��<M��<��<��<B��<���<֒�<"��<��<��<��<"��<֒�<���<B��<��<��<M��<A��<C��<:��<`   `   ��<)��<>��<)��<Q��<C��<9��<K��<	��<��<��<��<��<��<��<��<	��<K��<9��<C��<Q��<)��<>��<)��<`   `   Q��<g��<R��<7��<@��<��<��<H��<X��<7��<7��<@��<;��<@��<7��<7��<X��<H��<��<��<@��<7��<R��<g��<`   `   {��<P��<��<L��<G��<'��<i��<���<���<T��<���<ړ�<���<ړ�<���<T��<���<���<i��<'��<G��<L��<��<P��<`   `   b��<,��<��<f��<f��<���<��<ԓ�<���<���<ԓ�<���<���<���<ԓ�<���<���<ԓ�<��<���<f��<f��<��<,��<`   `   >��<5��<I��<i��<T��<���<���<o��<ӓ�<���<Г�<���<���<���<Г�<���<ӓ�<o��<���<���<T��<i��<I��<5��<`   `   0��<6��<M��<O��<I��<z��<���<���<
��<I��<	��<��<%��<��<	��<I��<
��<���<���<z��<I��<O��<M��<6��<`   `   7��<4��<3��<X��<���<���<��<'��<"��<`��<H��<w��<���<w��<H��<`��<"��<'��<��<���<���<X��<3��<4��<`   `   ?��<K��<,��<d��<ē�<���<ݓ�<��<��<^��<x��<���<���<���<x��<^��<��<��<ݓ�<���<ē�<d��<,��<K��<`   `   *��<R��<��<J��<ݓ�<���<���<*��<(��<���<ɔ�<���<���<���<ɔ�<���<(��<*��<���<���<ݓ�<J��<��<R��<`   `   ��<0��<��<?��<Γ�<œ�<��<���<k��<���<Ҕ�<���<���<���<Ҕ�<���<k��<���<��<œ�<Γ�<?��<��<0��<`   `   ���<>��<&��<I��<|��<���<��<!��<7��<N��<���<���<Ô�<���<���<N��<7��<!��<��<���<|��<I��<&��<>��<`   `   ��<<��<��<7��<M��<y��<�<ԓ�<>��<k��<���<���<���<���<���<k��<>��<ԓ�<�<y��<M��<7��<��<<��<`   `   ג�<��<͒�<��<7��<���<���<���<5��<���<���<���<���<���<���<���<5��<���<���<���<7��<��<͒�<��<`   `   Ԓ�<ݒ�<��<���<��<���<��<���<���<Z��<Z��<���<Ҕ�<���<Z��<Z��<���<���<��<���<��<���<��<ݒ�<`   `   ��<ޒ�<��<,��<��<+��<͓�<͓�<œ�<��<,��<b��<���<b��<,��<��<œ�<͓�<͓�<+��<��<,��<��<ޒ�<`   `   ��<���<���<���<��<��<���<��<˓�<��<T��<R��<&��<R��<T��<��<˓�<��<���<��<��<���<���<���<`   `   ���<}��<��<���<��<
��<K��<�<���<ߓ�<O��<8��<���<8��<O��<ߓ�<���<�<K��<
��<��<���<��<}��<`   `   M��<x��<���<���<���<0��<"��<F��<d��<���<�<��<-��<��<�<���<d��<F��<"��<0��<���<���<���<x��<`   `   Ñ�<%��<��<Y��<��<���<���<֑�<ؑ�<���<���<���<	��<���<���<���<ؑ�<֑�<���<���<��<Y��<��<%��<`   `   #��<	��<���<��<���<}��<S��<���<���<I��<��<���<���<���<��<I��<���<���<S��<}��<���<��<���<	��<`   `   ���<��<��<͐�<D��<p��<J��<���<���<���<֑�<��<ԑ�<��<֑�<���<���<���<J��<p��<D��<͐�<��<��<`   `   A��<`��<��<��<@��<2��<_��<���<���<��<���<x��<���<x��<���<��<���<���<_��<2��<@��<��<��<`��<`   `   m��<9��<��<@��<^��<1��<o��<{��<i��<���<~��<���<��<���<~��<���<i��<{��<o��<1��<^��<@��<��<9��<`   `   ,��<<��<Z��<���<y��<^��<���<���<{��<k��<���<���<Б�<���<���<k��<{��<���<���<^��<y��<���<Z��<<��<`   `   a��<���<���<���<p��<��<���<���<y��<j��<���<���<{��<���<���<j��<y��<���<���<��<p��<���<���<���<`   `   ���<���<~��<ȑ�<ґ�<���<���<���<���<���<���<^��<k��<^��<���<���<���<���<���<���<ґ�<ȑ�<~��<���<`   `   ���<�<���<��<Ց�<]��<���<Ñ�<���<���<���<g��<���<g��<���<���<���<Ñ�<���<]��<Ց�<��<���<�<`   `   ӑ�<��<��<��<���<n��<���<���<s��<���<���<e��<e��<e��<���<���<s��<���<���<n��<���<��<��<��<`   `   6��<\��<��<���<@��<��<���<ґ�<���<ב�<���<���<p��<���<���<ב�<���<ґ�<���<��<@��<���<��<\��<`   `   ���<���<C��<,��<9��<��<��<���<���<���<���<Ƒ�<���<Ƒ�<���<���<���<���<��<��<9��<,��<C��<���<`   `   {��<P��<X��<A��<��</��<��<��<͑�<���<���<u��<]��<u��<���<���<͑�<��<��</��<��<A��<X��<P��<`   `   i��<R��<w��<t��<W��<��<��<��<��<��<ё�<c��<���<c��<ё�<��<��<��<��<��<W��<t��<w��<R��<`   `   Ē�<���<w��<s��<E��<*��<��<��<���<���<Ƒ�<k��<đ�<k��<Ƒ�<���<���<��<��<*��<E��<s��<w��<���<`   `   ���<���<h��<���<R��<$��<C��<���<t��<���<���<[��<j��<[��<���<���<t��<���<C��<$��<R��<���<h��<���<`   `   x��<���<���<���<k��<!��<��<ɑ�<��<֑�<���<w��<U��<w��<���<֑�<��<ɑ�<��<!��<k��<���<���<���<`   `   ���<��<���<x��<l��<7��<��<Ց�<���<���<N��<>��<)��<>��<N��<���<���<Ց�<��<7��<l��<x��<���<��<`   `   `��<���<i��<k��<���<U��<*��<ɑ�<���<���<���<T��<B��<T��<���<���<���<ɑ�<*��<U��<���<k��<i��<���<`   `   W��<���<j��<���<���<���<���<���<���<���<p��<9��<8��<9��<p��<���<���<���<���<���<���<���<j��<���<`   `   |��<��<a��<\��<C��<Ց�<���<�<���<?��<���<��<ې�<��<���<?��<���<�<���<Ց�<C��<\��<a��<��<`   `   Z��</��<7��<��<��<��<���<���<^��<+��<a��<J��<���<J��<a��<+��<^��<���<���<��<��<��<7��</��<`   `   r��< ��<3��<��<���<ȑ�<|��<���<*��<`��<c��<��<��<��<c��<`��<*��<���<|��<ȑ�<���<��<3��< ��<`   `   |��<��<5��<��<���<Α�<~��<���<"��<���<��<Ԑ�<H��<Ԑ�<��<���<"��<���<~��<Α�<���<��<5��<��<`   `   	��<���<���<���<ؑ�<֑�<���<���<��<Y��<��<%��<Ñ�<%��<��<Y��<��<���<���<֑�<ؑ�<���<���<���<`   `   ���<���<��<I��<���<���<S��<}��<���<��<���<	��<#��<	��<���<��<���<}��<S��<���<���<I��<��<���<`   `   ԑ�<��<֑�<���<���<���<J��<p��<D��<͐�<��<��<���<��<��<͐�<D��<p��<J��<���<���<���<֑�<��<`   `   ���<x��<���<��<���<���<_��<2��<@��<��<��<`��<A��<`��<��<��<@��<2��<_��<���<���<��<���<x��<`   `   ��<���<~��<���<i��<{��<o��<1��<^��<@��<��<9��<m��<9��<��<@��<^��<1��<o��<{��<i��<���<~��<���<`   `   Б�<���<���<k��<{��<���<���<^��<y��<���<Z��<<��<+��<<��<Z��<���<y��<^��<���<���<{��<k��<���<���<`   `   {��<���<���<j��<y��<���<���<��<p��<���<���<���<a��<���<���<���<p��<��<���<���<y��<j��<���<���<`   `   k��<^��<���<���<���<���<���<���<ґ�<ȑ�<~��<���<���<���<~��<ȑ�<ґ�<���<���<���<���<���<���<^��<`   `   ���<g��<���<���<���<Ñ�<���<]��<Ց�<��<���<�<���<�<���<��<Ց�<]��<���<Ñ�<���<���<���<g��<`   `   e��<e��<���<���<s��<���<���<n��<���<��<��<��<ӑ�<��<��<��<���<n��<���<���<s��<���<���<e��<`   `   p��<���<���<ב�<���<ґ�<���<��<@��<���<��<\��<6��<\��<��<���<@��<��<���<ґ�<���<ב�<���<���<`   `   ���<Ƒ�<���<���<���<���<��<��<9��<,��<C��<���<���<���<C��<,��<9��<��<��<���<���<���<���<Ƒ�<`   `   ]��<u��<���<���<͑�<��<��</��<��<A��<X��<P��<{��<P��<X��<A��<��</��<��<��<͑�<���<���<u��<`   `   ���<c��<ё�<��<��<��<��<��<W��<t��<w��<R��<i��<R��<w��<t��<W��<��<��<��<��<��<ё�<c��<`   `   đ�<k��<Ƒ�<���<���<��<��<*��<E��<s��<w��<���<Ē�<���<w��<s��<E��<*��<��<��<���<���<Ƒ�<k��<`   `   j��<[��<���<���<t��<���<C��<$��<R��<���<h��<���<���<���<h��<���<R��<$��<C��<���<t��<���<���<[��<`   `   U��<w��<���<֑�<��<ɑ�<��<!��<k��<���<���<���<x��<���<���<���<k��<!��<��<ɑ�<��<֑�<���<w��<`   `   )��<>��<N��<���<���<Ց�<��<7��<l��<x��<���<��<���<��<���<x��<l��<7��<��<Ց�<���<���<N��<>��<`   `   B��<T��<���<���<���<ɑ�<*��<U��<���<k��<i��<���<`��<���<i��<k��<���<U��<*��<ɑ�<���<���<���<T��<`   `   8��<9��<p��<���<���<���<���<���<���<���<j��<���<W��<���<j��<���<���<���<���<���<���<���<p��<9��<`   `   ې�<��<���<?��<���<�<���<Ց�<C��<\��<a��<��<|��<��<a��<\��<C��<Ց�<���<�<���<?��<���<��<`   `   ���<J��<a��<+��<^��<���<���<��<��<��<7��</��<Z��</��<7��<��<��<��<���<���<^��<+��<a��<J��<`   `   ��<��<c��<`��<*��<���<|��<ȑ�<���<��<3��< ��<r��< ��<3��<��<���<ȑ�<|��<���<*��<`��<c��<��<`   `   H��<Ԑ�<��<���<"��<���<~��<Α�<���<��<5��<��<|��<��<5��<��<���<Α�<~��<���<"��<���<��<Ԑ�<`   `    ��<���<���<ҏ�<���<ˏ�<ߏ�<ˏ�<��<;��<���<E��<'��<E��<���<;��<��<ˏ�<ߏ�<ˏ�<���<ҏ�<���<���<`   `   I��<���<���<ȏ�<ݏ�<��<���<���<��<#��<��<��<��<��<��<#��<��<���<���<��<ݏ�<ȏ�<���<���<`   `   ���<���<���<���<��<���<ߏ�<���<��<��<���<��<��<��<���<��<��<���<ߏ�<���<��<���<���<���<`   `   X��<���<Տ�<��<��<���<��<���<���<��<	��<)��< ��<)��<	��<��<���<���<��<���<��<��<Տ�<���<`   `   ���<���<ˏ�<ڏ�<���<��<��<��<���<���<��<���<ȏ�<���<��<���<���<��<��<��<���<ڏ�<ˏ�<���<`   `   ��<���<���<��<ȏ�<؏�<��< ��<��<���<��<Ə�<���<Ə�<��<���<��< ��<��<؏�<ȏ�<��<���<���<`   `   ܏�<��<֏�<��<ɏ�<͏�<���<���<���<��<��<��<X��<��<��<��<���<���<���<͏�<ɏ�<��<֏�<��<`   `   	��<3��<���<ڏ�<���<��<��<܏�<��<��<ҏ�<�<3��<�<ҏ�<��<��<܏�<��<��<���<ڏ�<���<3��<`   `   (��<��<���<��<��<?��<��<"��<(��<��<��<���<��<���<��<��<(��<"��<��<?��<��<��<���<��<`   `   y��<��<+��<3��<��<O��<؏�<��<
��<�<��<@��<��<@��<��<�<
��<��<؏�<O��<��<3��<+��<��<`   `   o��<P��<k��<(��<[��<���<3��<��<$��<��<���<��<ȏ�<��<���<��<$��<��<3��<���<[��<(��<k��<P��<`   `   #��<B��<���<F��<F��<^��<=��<��<1��<#��<ҏ�<��<ۏ�<��<ҏ�<#��<1��<��<=��<^��<F��<F��<���<B��<`   `   q��<���<���<o��<=��<*��<��<��<���<���<��<��<��<��<��<���<���<��<��<*��<=��<o��<���<���<`   `   Ő�<א�<���<���<���<o��<K��<h��<��<��<��<؏�<"��<؏�<��<��<��<h��<K��<o��<���<���<���<א�<`   `   ���<ؐ�<���<���<���<L��<`��<���<��<��<���<���<:��<���<���<��<��<���<`��<L��<���<���<���<ؐ�<`   `   ���<ؐ�<���<���<���<A��<N��<I��<#��<��<��<���<��<���<��<��<#��<I��<N��<A��<���<���<���<ؐ�<`   `   ʐ�<֐�<���<ڐ�<���<���<F��<��<��<ʏ�<ҏ�<��<4��<��<ҏ�<ʏ�<��<��<F��<���<���<ڐ�<���<֐�<`   `   ֐�<���<���<���<X��<v��<F��<1��<���<���<ȏ�<ȏ�<��<ȏ�<ȏ�<���<���<1��<F��<v��<X��<���<���<���<`   `   Ӑ�<���<���<i��<!��<V��<��<��<��<Ǐ�<��<���<��<���<��<Ǐ�<��<��<��<V��<!��<i��<���<���<`   `   ���<���<���<O��<@��<���<��<���<���<�<ӏ�<͏�<��<͏�<ӏ�<�<���<���<��<���<@��<O��<���<���<`   `   ���<���<���<b��<Z��<u��<D��<��<��<���<���<���<���<���<���<���<��<��<D��<u��<Z��<b��<���<���<`   `   ���<���<|��<w��<S��<��<��<��<ŏ�<���<�<ˏ�<{��<ˏ�<�<���<ŏ�<��<��<��<S��<w��<|��<���<`   `   ���<N��<<��<"��<9��<���<��<���<���<���<`��<���<���<���<`��<���<���<���<��<���<9��<"��<<��<N��<`   `   T��<;��<v��<��<��<��<���<ʏ�<���<���<C��<���<s��<���<C��<���<���<ʏ�<���<��<��<��<v��<;��<`   `   '��<E��<���<;��<��<ˏ�<ߏ�<ˏ�<���<ҏ�<���<���< ��<���<���<ҏ�<���<ˏ�<ߏ�<ˏ�<��<;��<���<E��<`   `   ��<��<��<#��<��<���<���<��<ݏ�<ȏ�<���<���<I��<���<���<ȏ�<ݏ�<��<���<���<��<#��<��<��<`   `   ��<��<���<��<��<���<ߏ�<���<��<���<���<���<���<���<���<���<��<���<ߏ�<���<��<��<���<��<`   `    ��<)��<	��<��<���<���<��<���<��<��<Տ�<���<X��<���<Տ�<��<��<���<��<���<���<��<	��<)��<`   `   ȏ�<���<��<���<���<��<��<��<���<ڏ�<ˏ�<���<���<���<ˏ�<ڏ�<���<��<��<��<���<���<��<���<`   `   ���<Ə�<��<���<��< ��<��<؏�<ȏ�<��<���<���<��<���<���<��<ȏ�<؏�<��< ��<��<���<��<Ə�<`   `   X��<��<��<��<���<���<���<͏�<ɏ�<��<֏�<��<܏�<��<֏�<��<ɏ�<͏�<���<���<���<��<��<��<`   `   3��<�<ҏ�<��<��<܏�<��<��<���<ڏ�<���<3��<	��<3��<���<ڏ�<���<��<��<܏�<��<��<ҏ�<�<`   `   ��<���<��<��<(��<"��<��<?��<��<��<���<��<(��<��<���<��<��<?��<��<"��<(��<��<��<���<`   `   ��<@��<��<�<
��<��<؏�<O��<��<3��<+��<��<y��<��<+��<3��<��<O��<؏�<��<
��<�<��<@��<`   `   ȏ�<��<���<��<$��<��<3��<���<[��<(��<k��<P��<o��<P��<k��<(��<[��<���<3��<��<$��<��<���<��<`   `   ۏ�<��<ҏ�<#��<1��<��<=��<^��<F��<F��<���<B��<#��<B��<���<F��<F��<^��<=��<��<1��<#��<ҏ�<��<`   `   ��<��<��<���<���<��<��<*��<=��<o��<���<���<q��<���<���<o��<=��<*��<��<��<���<���<��<��<`   `   "��<؏�<��<��<��<h��<K��<o��<���<���<���<א�<Ő�<א�<���<���<���<o��<K��<h��<��<��<��<؏�<`   `   :��<���<���<��<��<���<`��<L��<���<���<���<ؐ�<���<ؐ�<���<���<���<L��<`��<���<��<��<���<���<`   `   ��<���<��<��<#��<I��<N��<A��<���<���<���<ؐ�<���<ؐ�<���<���<���<A��<N��<I��<#��<��<��<���<`   `   4��<��<ҏ�<ʏ�<��<��<F��<���<���<ڐ�<���<֐�<ʐ�<֐�<���<ڐ�<���<���<F��<��<��<ʏ�<ҏ�<��<`   `   ��<ȏ�<ȏ�<���<���<1��<F��<v��<X��<���<���<���<֐�<���<���<���<X��<v��<F��<1��<���<���<ȏ�<ȏ�<`   `   ��<���<��<Ǐ�<��<��<��<V��<!��<i��<���<���<Ӑ�<���<���<i��<!��<V��<��<��<��<Ǐ�<��<���<`   `   ��<͏�<ӏ�<�<���<���<��<���<@��<O��<���<���<���<���<���<O��<@��<���<��<���<���<�<ӏ�<͏�<`   `   ���<���<���<���<��<��<D��<u��<Z��<b��<���<���<���<���<���<b��<Z��<u��<D��<��<��<���<���<���<`   `   {��<ˏ�<�<���<ŏ�<��<��<��<S��<w��<|��<���<���<���<|��<w��<S��<��<��<��<ŏ�<���<�<ˏ�<`   `   ���<���<`��<���<���<���<��<���<9��<"��<<��<N��<���<N��<<��<"��<9��<���<��<���<���<���<`��<���<`   `   s��<���<C��<���<���<ʏ�<���<��<��<��<v��<;��<T��<;��<v��<��<��<��<���<ʏ�<���<���<C��<���<`   `   ���<E��<��<��<L��<��<J��<U��<���<p��<7��<���<���<���<7��<p��<���<U��<J��<��<L��<��<��<E��<`   `   ��<"��<���<!��<��<���<���<X��<���<���<m��<���<���<���<m��<���<���<X��<���<���<��<!��<���<"��<`   `   ���<��<��<$��<��<ݍ�<r��<m��<R��<o��<���<���<=��<���<���<o��<R��<m��<r��<ݍ�<��<$��<��<��<`   `   ��<֍�<��<	��<��<I��<B��<���<l��<.��<Y��<���<J��<���<Y��<.��<l��<���<B��<I��<��<	��<��<֍�<`   `   W��<C��<k��<��<���<V��<��<C��<���<3��<J��<���<i��<���<J��<3��<���<C��<��<V��<���<��<k��<C��<`   `   j��<T��<A��<��<8��<e��<&��<=��<_��<5��<S��<b��<3��<b��<S��<5��<_��<=��<&��<e��<8��<��<A��<T��<`   `   ��<%��<4��<z��<���<q��<|��<u��<Q��<K��<n��<_��<R��<_��<n��<K��<Q��<u��<|��<q��<���<z��<4��<%��<`   `   ��<w��<|��<i��<_��<B��<B��<E��<D��<T��<d��<E��<Z��<E��<d��<T��<D��<E��<B��<B��<_��<i��<|��<w��<`   `   ���<���<���<}��<u��<���<H��<@��<U��<M��<P��<!��<!��<!��<P��<M��<U��<@��<H��<���<u��<}��<���<���<`   `   ̎�<���<���<���<z��<���<l��<���<���<e��<_��<F��<@��<F��<_��<e��<���<���<l��<���<z��<���<���<���<`   `   ���<���<���<���<K��<��<f��<���<N��<q��<\��<Z��<\��<Z��<\��<q��<N��<���<f��<��<K��<���<���<���<`   `   ���<���<���<��<̎�<q��<���<f��<:��<���<i��<i��<M��<i��<i��<���<:��<f��<���<q��<̎�<��<���<���<`   `   <��<��<���<Վ�<��<���<Ҏ�<���<���<���<Q��<d��<-��<d��<Q��<���<���<���<Ҏ�<���<��<Վ�<���<��<`   `   ��<Ҏ�<���<���<���<���<���<g��<���<]��<8��<_��<+��<_��<8��<]��<���<g��<���<���<���<���<���<Ҏ�<`   `   ���<Ύ�<���<ێ�<���<͎�<���<&��<���<o��<a��<w��<;��<w��<a��<o��<���<&��<���<͎�<���<ێ�<���<Ύ�<`   `   ܎�<��<��<׎�<���<��<���<N��<���<c��<T��<_��<��<_��<T��<c��<���<N��<���<��<���<׎�<��<��<`   `   ��<���<��<���<���<֎�<���<}��<���<X��<e��<I��<���<I��<e��<X��<���<}��<���<֎�<���<���<��<���<`   `   ��<���<ގ�<���<ώ�<���<���<���<o��<���<���<8��<0��<8��<���<���<o��<���<���<���<ώ�<���<ގ�<���<`   `   ,��<ǎ�<��<N��<��<���<��<���<^��<l��<@��<��<)��<��<@��<l��<^��<���<��<���<��<N��<��<ǎ�<`   `   #��<���<Ȏ�< ��<���<���<���<���<W��<-��<��<��<��<��<��<-��<W��<���<���<���<���< ��<Ȏ�<���<`   `   ���<���<���<���<���<���<���<)��<:��<k��<]��<6��<4��<6��<]��<k��<:��<)��<���<���<���<���<���<���<`   `   ���<َ�<���<ǎ�<���<r��<y��<��<3��<���<
��<���<
��<���<
��<���<3��<��<y��<r��<���<ǎ�<���<َ�<`   `   ���<܎�<֎�<���<���<���<���<3��<v��<\��<��<��<���<��<��<\��<v��<3��<���<���<���<���<֎�<܎�<`   `   ���<���<{��<f��<���<���<T��<)��<l��<��<>��<���<���<���<>��<��<l��<)��<T��<���<���<f��<{��<���<`   `   ���<���<7��<p��<���<U��<J��<��<L��<��<��<E��<���<E��<��<��<L��<��<J��<U��<���<p��<7��<���<`   `   ���<���<m��<���<���<X��<���<���<��<!��<���<"��<��<"��<���<!��<��<���<���<X��<���<���<m��<���<`   `   =��<���<���<o��<R��<m��<r��<ݍ�<��<$��<��<��<���<��<��<$��<��<ݍ�<r��<m��<R��<o��<���<���<`   `   J��<���<Y��<.��<l��<���<B��<I��<��<	��<��<֍�<��<֍�<��<	��<��<I��<B��<���<l��<.��<Y��<���<`   `   i��<���<J��<3��<���<C��<��<V��<���<��<k��<C��<W��<C��<k��<��<���<V��<��<C��<���<3��<J��<���<`   `   3��<b��<S��<5��<_��<=��<&��<e��<8��<��<A��<T��<j��<T��<A��<��<8��<e��<&��<=��<_��<5��<S��<b��<`   `   R��<_��<n��<K��<Q��<u��<|��<q��<���<z��<4��<%��<��<%��<4��<z��<���<q��<|��<u��<Q��<K��<n��<_��<`   `   Z��<E��<d��<T��<D��<E��<B��<B��<_��<i��<|��<w��<��<w��<|��<i��<_��<B��<B��<E��<D��<T��<d��<E��<`   `   !��<!��<P��<M��<U��<@��<H��<���<u��<}��<���<���<���<���<���<}��<u��<���<H��<@��<U��<M��<P��<!��<`   `   @��<F��<_��<e��<���<���<l��<���<z��<���<���<���<̎�<���<���<���<z��<���<l��<���<���<e��<_��<F��<`   `   \��<Z��<\��<q��<N��<���<f��<��<K��<���<���<���<���<���<���<���<K��<��<f��<���<N��<q��<\��<Z��<`   `   M��<i��<i��<���<:��<f��<���<q��<̎�<��<���<���<���<���<���<��<̎�<q��<���<f��<:��<���<i��<i��<`   `   -��<d��<Q��<���<���<���<Ҏ�<���<��<Վ�<���<��<<��<��<���<Վ�<��<���<Ҏ�<���<���<���<Q��<d��<`   `   +��<_��<8��<]��<���<g��<���<���<���<���<���<Ҏ�<��<Ҏ�<���<���<���<���<���<g��<���<]��<8��<_��<`   `   ;��<w��<a��<o��<���<&��<���<͎�<���<ێ�<���<Ύ�<���<Ύ�<���<ێ�<���<͎�<���<&��<���<o��<a��<w��<`   `   ��<_��<T��<c��<���<N��<���<��<���<׎�<��<��<܎�<��<��<׎�<���<��<���<N��<���<c��<T��<_��<`   `   ���<I��<e��<X��<���<}��<���<֎�<���<���<��<���<��<���<��<���<���<֎�<���<}��<���<X��<e��<I��<`   `   0��<8��<���<���<o��<���<���<���<ώ�<���<ގ�<���<��<���<ގ�<���<ώ�<���<���<���<o��<���<���<8��<`   `   )��<��<@��<l��<^��<���<��<���<��<N��<��<ǎ�<,��<ǎ�<��<N��<��<���<��<���<^��<l��<@��<��<`   `   ��<��<��<-��<W��<���<���<���<���< ��<Ȏ�<���<#��<���<Ȏ�< ��<���<���<���<���<W��<-��<��<��<`   `   4��<6��<]��<k��<:��<)��<���<���<���<���<���<���<���<���<���<���<���<���<���<)��<:��<k��<]��<6��<`   `   
��<���<
��<���<3��<��<y��<r��<���<ǎ�<���<َ�<���<َ�<���<ǎ�<���<r��<y��<��<3��<���<
��<���<`   `   ���<��<��<\��<v��<3��<���<���<���<���<֎�<܎�<���<܎�<֎�<���<���<���<���<3��<v��<\��<��<��<`   `   ���<���<>��<��<l��<)��<T��<���<���<f��<{��<���<���<���<{��<f��<���<���<T��<)��<l��<��<>��<���<`   `   ���<p��<g��<���<���<���<Ռ�<��<ڌ�<��<��<���<��<���<��<��<ڌ�<��<Ռ�<���<���<���<g��<p��<`   `   ���<o��<���<���<ƌ�<��<���<Č�<���<���<���<���<ٌ�<���<���<���<���<Č�<���<��<ƌ�<���<���<o��<`   `   m��<t��<��<���<���<���<���<���<���<Ɍ�<��<��<ٌ�<��<��<Ɍ�<���<���<���<���<���<���<��<t��<`   `   Ќ�<���<���<���<��<���<���<ی�<ь�<��<���<���<���<���<���<��<ь�<ی�<���<���<��<���<���<���<`   `   ���<���<���<ߌ�<��<���<���<Ԍ�<Ԍ�<��<Ō�<���<��<���<Ō�<��<Ԍ�<Ԍ�<���<���<��<ߌ�<���<���<`   `   ���<���<Ì�<֌�<���<���<��<���<���<��<ь�<��<���<��<ь�<��<���<���<��<���<���<֌�<Ì�<���<`   `   ��<���<���<Ì�<���<���<���<��<���<���<���<���<~��<���<���<���<���<��<���<���<���<Ì�<���<���<`   `   ��<���<���<Ȍ�<֌�<���<ό�<��<��<ތ�<܌�<��<Ȍ�<��<܌�<ތ�<��<��<ό�<���<֌�<Ȍ�<���<���<`   `   ���<ʌ�<���<���<��<���<ڌ�<ǌ�<���<Ԍ�<���<��<��<��<���<Ԍ�<���<ǌ�<ڌ�<���<��<���<���<ʌ�<`   `   Ό�<��<ߌ�<݌�<��<���<��<���<���<���<���<���<��<���<���<���<���<���<��<���<��<݌�<ߌ�<��<`   `   ��<#��<���<��</��<��< ��<���<���<��<��<ˌ�<���<ˌ�<��<��<���<���< ��<��</��<��<���<#��<`   `   ��<D��<��<׌�<#��<��<���<��<���<���<���<Ό�<ˌ�<Ό�<���<���<���<��<���<��<#��<׌�<��<D��<`   `   ٌ�<��<.��<
��<��<���<��<��<���<���<���<܌�<ˌ�<܌�<���<���<���<��<��<���<��<
��<.��<��<`   `   ��<(��<N��<B��<���<��<��<��<��<ی�<׌�<��<���<��<׌�<ی�<��<��<��<��<���<B��<N��<(��<`   `   ���<O��<5��<G��<#��<��<;��<���<ӌ�<Ō�<ڌ�<��<���<��<ڌ�<Ō�<ӌ�<���<;��<��<#��<G��<5��<O��<`   `   ��<��<��<@��<5��<��<#��<+��<ٌ�<���<���<��<�<��<���<���<ٌ�<+��<#��<��<5��<@��<��<��<`   `   M��<4��<O��<8��<:��<̌�<���<��<���<���<���<ό�<���<ό�<���<���<���<��<���<̌�<:��<8��<O��<4��<`   `   F��<s��<`��<��<H��<��<���<Ό�<���<��<���<���<ی�<���<���<��<���<Ό�<���<��<H��<��<`��<s��<`   `    ��<E��<��<���<#��< ��<���<���<���<̌�<���<���<(��<���<���<̌�<���<���<���< ��<#��<���<��<E��<`   `   )��<;��<'��<��<��<��<Ҍ�<ʌ�<Ҍ�<���<͌�<݌�<���<݌�<͌�<���<Ҍ�<ʌ�<Ҍ�<��<��<��<'��<;��<`   `   J��<_��<E��<J��<4��<��<Ɍ�<��<���<���<���<���<���<���<���<���<���<��<Ɍ�<��<4��<J��<E��<_��<`   `   ��<3��<��<��<���<��<��<#��<���<P��<���<���<��<���<���<P��<���<#��<��<��<���<��<��<3��<`   `   ��<��<��<��<���<���<ό�<��<���<���<Ҍ�<q��<���<q��<Ҍ�<���<���<��<ό�<���<���<��<��<��<`   `   ��<��<(��<C��<Ќ�<���<���<���<���<���<Ō�<Z��<}��<Z��<Ō�<���<���<���<���<���<Ќ�<C��<(��<��<`   `   ��<���<��<��<ڌ�<��<Ռ�<���<���<���<g��<p��<���<p��<g��<���<���<���<Ռ�<��<ڌ�<��<��<���<`   `   ٌ�<���<���<���<���<Č�<���<��<ƌ�<���<���<o��<���<o��<���<���<ƌ�<��<���<Č�<���<���<���<���<`   `   ٌ�<��<��<Ɍ�<���<���<���<���<���<���<��<t��<m��<t��<��<���<���<���<���<���<���<Ɍ�<��<��<`   `   ���<���<���<��<ь�<ی�<���<���<��<���<���<���<Ќ�<���<���<���<��<���<���<ی�<ь�<��<���<���<`   `   ��<���<Ō�<��<Ԍ�<Ԍ�<���<���<��<ߌ�<���<���<���<���<���<ߌ�<��<���<���<Ԍ�<Ԍ�<��<Ō�<���<`   `   ���<��<ь�<��<���<���<��<���<���<֌�<Ì�<���<���<���<Ì�<֌�<���<���<��<���<���<��<ь�<��<`   `   ~��<���<���<���<���<��<���<���<���<Ì�<���<���<��<���<���<Ì�<���<���<���<��<���<���<���<���<`   `   Ȍ�<��<܌�<ތ�<��<��<ό�<���<֌�<Ȍ�<���<���<��<���<���<Ȍ�<֌�<���<ό�<��<��<ތ�<܌�<��<`   `   ��<��<���<Ԍ�<���<ǌ�<ڌ�<���<��<���<���<ʌ�<���<ʌ�<���<���<��<���<ڌ�<ǌ�<���<Ԍ�<���<��<`   `   ��<���<���<���<���<���<��<���<��<݌�<ߌ�<��<Ό�<��<ߌ�<݌�<��<���<��<���<���<���<���<���<`   `   ���<ˌ�<��<��<���<���< ��<��</��<��<���<#��<��<#��<���<��</��<��< ��<���<���<��<��<ˌ�<`   `   ˌ�<Ό�<���<���<���<��<���<��<#��<׌�<��<D��<��<D��<��<׌�<#��<��<���<��<���<���<���<Ό�<`   `   ˌ�<܌�<���<���<���<��<��<���<��<
��<.��<��<ٌ�<��<.��<
��<��<���<��<��<���<���<���<܌�<`   `   ���<��<׌�<ی�<��<��<��<��<���<B��<N��<(��<��<(��<N��<B��<���<��<��<��<��<ی�<׌�<��<`   `   ���<��<ڌ�<Ō�<ӌ�<���<;��<��<#��<G��<5��<O��<���<O��<5��<G��<#��<��<;��<���<ӌ�<Ō�<ڌ�<��<`   `   �<��<���<���<ٌ�<+��<#��<��<5��<@��<��<��<��<��<��<@��<5��<��<#��<+��<ٌ�<���<���<��<`   `   ���<ό�<���<���<���<��<���<̌�<:��<8��<O��<4��<M��<4��<O��<8��<:��<̌�<���<��<���<���<���<ό�<`   `   ی�<���<���<��<���<Ό�<���<��<H��<��<`��<s��<F��<s��<`��<��<H��<��<���<Ό�<���<��<���<���<`   `   (��<���<���<̌�<���<���<���< ��<#��<���<��<E��< ��<E��<��<���<#��< ��<���<���<���<̌�<���<���<`   `   ���<݌�<͌�<���<Ҍ�<ʌ�<Ҍ�<��<��<��<'��<;��<)��<;��<'��<��<��<��<Ҍ�<ʌ�<Ҍ�<���<͌�<݌�<`   `   ���<���<���<���<���<��<Ɍ�<��<4��<J��<E��<_��<J��<_��<E��<J��<4��<��<Ɍ�<��<���<���<���<���<`   `   ��<���<���<P��<���<#��<��<��<���<��<��<3��<��<3��<��<��<���<��<��<#��<���<P��<���<���<`   `   ���<q��<Ҍ�<���<���<��<ό�<���<���<��<��<��<��<��<��<��<���<���<ό�<��<���<���<Ҍ�<q��<`   `   }��<Z��<Ō�<���<���<���<���<���<Ќ�<C��<(��<��<��<��<(��<C��<Ќ�<���<���<���<���<���<Ō�<Z��<`   `   ���<��<,��<N��<��<#��<2��<g��<>��<Y��<���<{��<L��<{��<���<Y��<>��<g��<2��<#��<��<N��<,��<��<`   `   '��<��<U��<!��<��<(��<	��<z��<���<b��<T��<@��<B��<@��<T��<b��<���<z��<	��<(��<��<!��<U��<��<`   `   ˊ�<��<C��<���<��<H��<9��<~��<���<t��<5��<O��<���<O��<5��<t��<���<~��<9��<H��<��<���<C��<��<`   `   h��<p��<��<��<���<���<J��<D��<��<B��<]��<k��<���<k��<]��<B��<��<D��<J��<���<���<��<��<p��<`   `   <��<9��<��<O��<2��<���<���<b��<���<5��<`��<>��<4��<>��<`��<5��<���<b��<���<���<2��<O��<��<9��<`   `   %��<9��<>��<-��<9��<S��<h��<Q��<g��<g��<B��<R��<P��<R��<B��<g��<g��<Q��<h��<S��<9��<-��<>��<9��<`   `   X��<F��<[��<��<5��<t��<���<��<g��<X��<��<X��<T��<X��<��<X��<g��<��<���<t��<5��<��<[��<F��<`   `   ,��<��<g��<o��<���<���<S��<��<K��<?��<2��<U��<��<U��<2��<?��<K��<��<S��<���<���<o��<g��<��<`   `   {��<z��<���<u��<P��<a��<���<`��<\��<P��<H��<W��<��<W��<H��<P��<\��<`��<���<a��<P��<u��<���<z��<`   `   ���<���<���<h��<@��<,��<;��<+��<`��<I��<A��<O��<.��<O��<A��<I��<`��<+��<;��<,��<@��<h��<���<���<`   `   J��<m��<t��<���<��<���<A��<A��<���<A��<Q��<T��<@��<T��<Q��<A��<���<A��<A��<���<��<���<t��<m��<`   `   d��<|��<���<v��<:��<���<S��<p��<���<R��<\��<1��<1��<1��<\��<R��<���<p��<S��<���<:��<v��<���<|��<`   `   ���<���<���<���<_��<x��<L��<U��<K��<]��<z��<?��<i��<?��<z��<]��<K��<U��<L��<x��<_��<���<���<���<`   `   ���<���<���<���<�<���<q��<}��<)��<c��<d��<6��<���<6��<d��<c��<)��<}��<q��<���<�<���<���<���<`   `   ���<���<���<S��<���<k��<R��<���<P��<���<"��<��<N��<��<"��<���<P��<���<R��<k��<���<S��<���<���<`   `   ���<u��<���<q��<���<j��<A��<T��<M��<���<F��<&��<o��<&��<F��<���<M��<T��<A��<j��<���<q��<���<u��<`   `   ���<y��<���<���<���<���<���<b��<L��<���<d��<^��<T��<^��<d��<���<L��<b��<���<���<���<���<���<y��<`   `   ���<���<���<���<���<_��<���<{��<w��<\��<,��<@��<Ҋ�<@��<,��<\��<w��<{��<���<_��<���<���<���<���<`   `   w��<���<���<���<���<[��<���<t��<���<M��<$��<L��<���<L��<$��<M��<���<t��<���<[��<���<���<���<���<`   `   l��<���<���<���<p��<u��<���<=��<L��<M��<:��<E��<��<E��<:��<M��<L��<=��<���<u��<p��<���<���<���<`   `   \��<t��<���<z��<`��<���<[��<(��<9��<D��<-��<��<���<��<-��<D��<9��<(��<[��<���<`��<z��<���<t��<`   `   ���<���<���<{��<t��<���<,��<D��<T��<C��<^��<%��<Z��<%��<^��<C��<T��<D��<,��<���<t��<{��<���<���<`   `   ���<z��<Y��<���<z��<���<*��<B��<8��<<��<r��<��<b��<��<r��<<��<8��<B��<*��<���<z��<���<Y��<z��<`   `   |��<m��<U��<u��<R��<��<^��<P��<8��<O��<(��<Ɗ�<G��<Ɗ�<(��<O��<8��<P��<^��<��<R��<u��<U��<m��<`   `   L��<{��<���<Y��<>��<g��<2��<#��<��<N��<,��<��<���<��<,��<N��<��<#��<2��<g��<>��<Y��<���<{��<`   `   B��<@��<T��<b��<���<z��<	��<(��<��<!��<U��<��<'��<��<U��<!��<��<(��<	��<z��<���<b��<T��<@��<`   `   ���<O��<5��<t��<���<~��<9��<H��<��<���<C��<��<ˊ�<��<C��<���<��<H��<9��<~��<���<t��<5��<O��<`   `   ���<k��<]��<B��<��<D��<J��<���<���<��<��<p��<h��<p��<��<��<���<���<J��<D��<��<B��<]��<k��<`   `   4��<>��<`��<5��<���<b��<���<���<2��<O��<��<9��<<��<9��<��<O��<2��<���<���<b��<���<5��<`��<>��<`   `   P��<R��<B��<g��<g��<Q��<h��<S��<9��<-��<>��<9��<%��<9��<>��<-��<9��<S��<h��<Q��<g��<g��<B��<R��<`   `   T��<X��<��<X��<g��<��<���<t��<5��<��<[��<F��<X��<F��<[��<��<5��<t��<���<��<g��<X��<��<X��<`   `   ��<U��<2��<?��<K��<��<S��<���<���<o��<g��<��<,��<��<g��<o��<���<���<S��<��<K��<?��<2��<U��<`   `   ��<W��<H��<P��<\��<`��<���<a��<P��<u��<���<z��<{��<z��<���<u��<P��<a��<���<`��<\��<P��<H��<W��<`   `   .��<O��<A��<I��<`��<+��<;��<,��<@��<h��<���<���<���<���<���<h��<@��<,��<;��<+��<`��<I��<A��<O��<`   `   @��<T��<Q��<A��<���<A��<A��<���<��<���<t��<m��<J��<m��<t��<���<��<���<A��<A��<���<A��<Q��<T��<`   `   1��<1��<\��<R��<���<p��<S��<���<:��<v��<���<|��<d��<|��<���<v��<:��<���<S��<p��<���<R��<\��<1��<`   `   i��<?��<z��<]��<K��<U��<L��<x��<_��<���<���<���<���<���<���<���<_��<x��<L��<U��<K��<]��<z��<?��<`   `   ���<6��<d��<c��<)��<}��<q��<���<�<���<���<���<���<���<���<���<�<���<q��<}��<)��<c��<d��<6��<`   `   N��<��<"��<���<P��<���<R��<k��<���<S��<���<���<���<���<���<S��<���<k��<R��<���<P��<���<"��<��<`   `   o��<&��<F��<���<M��<T��<A��<j��<���<q��<���<u��<���<u��<���<q��<���<j��<A��<T��<M��<���<F��<&��<`   `   T��<^��<d��<���<L��<b��<���<���<���<���<���<y��<���<y��<���<���<���<���<���<b��<L��<���<d��<^��<`   `   Ҋ�<@��<,��<\��<w��<{��<���<_��<���<���<���<���<���<���<���<���<���<_��<���<{��<w��<\��<,��<@��<`   `   ���<L��<$��<M��<���<t��<���<[��<���<���<���<���<w��<���<���<���<���<[��<���<t��<���<M��<$��<L��<`   `   ��<E��<:��<M��<L��<=��<���<u��<p��<���<���<���<l��<���<���<���<p��<u��<���<=��<L��<M��<:��<E��<`   `   ���<��<-��<D��<9��<(��<[��<���<`��<z��<���<t��<\��<t��<���<z��<`��<���<[��<(��<9��<D��<-��<��<`   `   Z��<%��<^��<C��<T��<D��<,��<���<t��<{��<���<���<���<���<���<{��<t��<���<,��<D��<T��<C��<^��<%��<`   `   b��<��<r��<<��<8��<B��<*��<���<z��<���<Y��<z��<���<z��<Y��<���<z��<���<*��<B��<8��<<��<r��<��<`   `   G��<Ɗ�<(��<O��<8��<P��<^��<��<R��<u��<U��<m��<|��<m��<U��<u��<R��<��<^��<P��<8��<O��<(��<Ɗ�<`   `   Q��<҉�<��<���<׉�<͉�<��<���<ԉ�<��<��<"��<��<"��<��<��<ԉ�<���<��<͉�<׉�<���<��<҉�<`   `   ���<Չ�<���<���<ى�<ˉ�<��<���<���<݉�<���<���<��<���<���<݉�<���<���<��<ˉ�<ى�<���<���<Չ�<`   `   މ�<׉�<q��<���<��<���<��<���<���<Ɖ�<؉�<���<���<���<؉�<Ɖ�<���<���<��<���<��<���<q��<׉�<`   `   n��<���<���<��<���<щ�<܉�<���<��<׉�<
��<��<���<��<
��<׉�<��<���<܉�<щ�<���<��<���<���<`   `   w��<ى�<���<É�<ۉ�<���<���<���<��<���<��<��<���<��<��<���<��<���<���<���<ۉ�<É�<���<ى�<`   `   ��<���<��<ʉ�<���<���<���<��<��<���<ԉ�<߉�<ŉ�<߉�<ԉ�<���<��<��<���<���<���<ʉ�<��<���<`   `   ܉�<���<��<ۉ�<���<ŉ�<�<��<ԉ�<ԉ�<���<��<��<��<���<ԉ�<ԉ�<��<�<ŉ�<���<ۉ�<��<���<`   `   ���<���<��<։�<���<���<Ӊ�<��<���<Љ�<��<ɉ�<҉�<ɉ�<��<Љ�<���<��<Ӊ�<���<���<։�<��<���<`   `   ��<��<ԉ�<Љ�<։�<���<ǉ�<��<��<��<��<։�<���<։�<��<��<��<��<ǉ�<���<։�<Љ�<ԉ�<��<`   `   ĉ�<Љ�<���<��<��<���<���<��<��<ɉ�<��<��<ˉ�<��<��<ɉ�<��<��<���<���<��<��<���<Љ�<`   `   ��<��<։�<#��<؉�<��<��<Ӊ�<ɉ�<���<��<��<��<��<��<���<ɉ�<Ӊ�<��<��<؉�<#��<։�<��<`   `   T��<��<��<C��<։�<���<
��<��<ω�<ˉ�<��<Ή�<��<Ή�<��<ˉ�<ω�<��<
��<���<։�<C��<��<��<`   `   ^��<��<Ӊ�<$��<��<��<��<��<͉�<ۉ�<߉�<���<܉�<���<߉�<ۉ�<͉�<��<��<��<��<$��<Ӊ�<��<`   `   ��<��<ډ�<��<���<���<���<��<���<ω�<݉�<ω�<��<ω�<݉�<ω�<���<��<���<���<���<��<ډ�<��<`   `   ���<��<B��<��<���<���<׉�<���<��<���<��<��<
��<��<��<���<��<���<׉�<���<���<��<B��<��<`   `   ��<M��<{��<��<���<F��<���<ۉ�<̉�<���<Љ�<ȉ�<ȉ�<ȉ�<Љ�<���<̉�<ۉ�<���<F��<���<��<{��<M��<`   `   t��<*��<���<؉�<ȉ�<A��<��<���<ډ�<���<�<���<Љ�<���<�<���<ډ�<���<��<A��<ȉ�<؉�<���<*��<`   `   =��<ډ�<͉�<��<ى�<��<ˉ�<ȉ�<͉�<���<���<��<���<��<���<���<͉�<ȉ�<ˉ�<��<ى�<��<͉�<ډ�<`   `   C��<��<��<d��<1��<��<ĉ�<ȉ�<ۉ�<ŉ�<��<މ�<���<މ�<��<ŉ�<ۉ�<ȉ�<ĉ�<��<1��<d��<��<��<`   `   ���<&��<��<��<)��<��<���<��<ȉ�<։�<���<މ�<5��<މ�<���<։�<ȉ�<��<���<��<)��<��<��<&��<`   `   @��<��<ˉ�<��<ډ�<ȉ�<���<��<���<��<���<Ή�<4��<Ή�<���<��<���<��<���<ȉ�<ډ�<��<ˉ�<��<`   `   ��<���<5��<!��<ĉ�<҉�<��<ԉ�<މ�<��<���<���<o��<���<���<��<މ�<ԉ�<��<҉�<ĉ�<!��<5��<���<`   `   ���<��<&��<��<݉�<ԉ�<͉�<���<��<��<���<ԉ�<���<ԉ�<���<��<��<���<͉�<ԉ�<݉�<��<&��<��<`   `   ͉�<��<���<ԉ�<���<щ�<��<��<��<���<���<���<���<���<���<���<��<��<��<щ�<���<ԉ�<���<��<`   `   ��<"��<��<��<ԉ�<���<��<͉�<׉�<���<��<҉�<Q��<҉�<��<���<׉�<͉�<��<���<ԉ�<��<��<"��<`   `   ��<���<���<݉�<���<���<��<ˉ�<ى�<���<���<Չ�<���<Չ�<���<���<ى�<ˉ�<��<���<���<݉�<���<���<`   `   ���<���<؉�<Ɖ�<���<���<��<���<��<���<q��<׉�<މ�<׉�<q��<���<��<���<��<���<���<Ɖ�<؉�<���<`   `   ���<��<
��<׉�<��<���<܉�<щ�<���<��<���<���<n��<���<���<��<���<щ�<܉�<���<��<׉�<
��<��<`   `   ���<��<��<���<��<���<���<���<ۉ�<É�<���<ى�<w��<ى�<���<É�<ۉ�<���<���<���<��<���<��<��<`   `   ŉ�<߉�<ԉ�<���<��<��<���<���<���<ʉ�<��<���<��<���<��<ʉ�<���<���<���<��<��<���<ԉ�<߉�<`   `   ��<��<���<ԉ�<ԉ�<��<�<ŉ�<���<ۉ�<��<���<܉�<���<��<ۉ�<���<ŉ�<�<��<ԉ�<ԉ�<���<��<`   `   ҉�<ɉ�<��<Љ�<���<��<Ӊ�<���<���<։�<��<���<���<���<��<։�<���<���<Ӊ�<��<���<Љ�<��<ɉ�<`   `   ���<։�<��<��<��<��<ǉ�<���<։�<Љ�<ԉ�<��<��<��<ԉ�<Љ�<։�<���<ǉ�<��<��<��<��<։�<`   `   ˉ�<��<��<ɉ�<��<��<���<���<��<��<���<Љ�<ĉ�<Љ�<���<��<��<���<���<��<��<ɉ�<��<��<`   `   ��<��<��<���<ɉ�<Ӊ�<��<��<؉�<#��<։�<��<��<��<։�<#��<؉�<��<��<Ӊ�<ɉ�<���<��<��<`   `   ��<Ή�<��<ˉ�<ω�<��<
��<���<։�<C��<��<��<T��<��<��<C��<։�<���<
��<��<ω�<ˉ�<��<Ή�<`   `   ܉�<���<߉�<ۉ�<͉�<��<��<��<��<$��<Ӊ�<��<^��<��<Ӊ�<$��<��<��<��<��<͉�<ۉ�<߉�<���<`   `   ��<ω�<݉�<ω�<���<��<���<���<���<��<ډ�<��<��<��<ډ�<��<���<���<���<��<���<ω�<݉�<ω�<`   `   
��<��<��<���<��<���<׉�<���<���<��<B��<��<���<��<B��<��<���<���<׉�<���<��<���<��<��<`   `   ȉ�<ȉ�<Љ�<���<̉�<ۉ�<���<F��<���<��<{��<M��<��<M��<{��<��<���<F��<���<ۉ�<̉�<���<Љ�<ȉ�<`   `   Љ�<���<�<���<ډ�<���<��<A��<ȉ�<؉�<���<*��<t��<*��<���<؉�<ȉ�<A��<��<���<ډ�<���<�<���<`   `   ���<��<���<���<͉�<ȉ�<ˉ�<��<ى�<��<͉�<ډ�<=��<ډ�<͉�<��<ى�<��<ˉ�<ȉ�<͉�<���<���<��<`   `   ���<މ�<��<ŉ�<ۉ�<ȉ�<ĉ�<��<1��<d��<��<��<C��<��<��<d��<1��<��<ĉ�<ȉ�<ۉ�<ŉ�<��<މ�<`   `   5��<މ�<���<։�<ȉ�<��<���<��<)��<��<��<&��<���<&��<��<��<)��<��<���<��<ȉ�<։�<���<މ�<`   `   4��<Ή�<���<��<���<��<���<ȉ�<ډ�<��<ˉ�<��<@��<��<ˉ�<��<ډ�<ȉ�<���<��<���<��<���<Ή�<`   `   o��<���<���<��<މ�<ԉ�<��<҉�<ĉ�<!��<5��<���<��<���<5��<!��<ĉ�<҉�<��<ԉ�<މ�<��<���<���<`   `   ���<ԉ�<���<��<��<���<͉�<ԉ�<݉�<��<&��<��<���<��<&��<��<݉�<ԉ�<͉�<���<��<��<���<ԉ�<`   `   ���<���<���<���<��<��<��<щ�<���<ԉ�<���<��<͉�<��<���<ԉ�<���<щ�<��<��<��<���<���<���<`   `   ��<N��<j��<s��<c��<_��<���<���<Έ�<���<g��<b��<P��<b��<g��<���<Έ�<���<���<_��<c��<s��<j��<N��<`   `   T��<p��<R��<^��<[��<?��<r��<���<���<���<���<q��<���<q��<���<���<���<���<r��<?��<[��<^��<R��<p��<`   `   ��<y��<Z��<s��<*��<��<C��<s��<c��<Z��<���<x��<���<x��<���<Z��<c��<s��<C��<��<*��<s��<Z��<y��<`   `   7��<i��<|��<a��<��<p��<w��<r��<���<g��<j��<t��<���<t��<j��<g��<���<r��<w��<p��<��<a��<|��<i��<`   `   _��<���<]��<5��<.��<���<���<Y��<���<s��<Y��<|��<Ĉ�<|��<Y��<s��<���<Y��<���<���<.��<5��<]��<���<`   `   n��<W��<D��<o��<]��<;��<X��<B��<��<q��<~��<V��<���<V��<~��<q��<��<B��<X��<;��<]��<o��<D��<W��<`   `   u��<@��<W��<���<{��<`��<���<���<"��<���<���<-��<\��<-��<���<���<"��<���<���<`��<{��<���<W��<@��<`   `   Έ�<���<|��<c��<���<���<{��<���<g��<���<X��<S��<���<S��<X��<���<g��<���<{��<���<���<c��<|��<���<`   `   b��<���<���<r��<���<���<8��<E��<e��<t��<O��<���<���<���<O��<t��<e��<E��<8��<���<���<r��<���<���<`   `   :��<���<���<���<���<���<���<~��<n��<���<j��<Z��<~��<Z��<j��<���<n��<~��<���<���<���<���<���<���<`   `   ���<و�<���<\��<g��<f��<j��<u��<y��<���<z��<4��<W��<4��<z��<���<y��<u��<j��<f��<g��<\��<���<و�<`   `   $��<���<���<c��<���<}��<R��<���<���<���<w��<c��<���<c��<w��<���<���<���<R��<}��<���<c��<���<���<`   `   ��<���<���<���<���<���<p��<w��<���<s��<f��<���<���<���<f��<s��<���<w��<p��<���<���<���<���<���<`   `   ���<Ɉ�<Ĉ�<���<`��<e��<���<E��<���<|��<W��<o��<��<o��<W��<|��<���<E��<���<e��<`��<���<Ĉ�<Ɉ�<`   `   ��<���<Y��<ƈ�<���<���<È�<d��<���<c��<���<���<��<���<���<c��<���<d��<È�<���<���<ƈ�<Y��<���<`   `   ���<x��<,��<���<���<W��<��<���<���<g��<���<���<G��<���<���<g��<���<���<��<W��<���<���<,��<x��<`   `   H��<���<���<ш�<���<M��<E��<���<���<���<w��<&��<{��<&��<w��<���<���<���<E��<M��<���<ш�<���<���<`   `   ���<���<؈�<���<���<���<���<���<���<}��<q��<8��<ˈ�<8��<q��<}��<���<���<���<���<���<���<؈�<���<`   `   Q��<���<���<2��<>��<͈�<���<��<j��<z��<{��<��<c��<��<{��<z��<j��<��<���<͈�<>��<2��<���<���<`   `   /��<���<���<O��<y��<���<Q��<���<���<���<l��<��<-��<��<l��<���<���<���<Q��<���<y��<O��<���<���<`   `   ���<���<͈�<���<��<���<R��<���<W��<Q��<q��<y��<T��<y��<q��<Q��<W��<���<R��<���<��<���<͈�<���<`   `   ���<j��<_��<h��<���<���<���<���<U��<b��<v��<���<��<���<v��<b��<U��<���<���<���<���<h��<_��<j��<`   `   ���<���<~��<R��<s��<b��<���<J��<e��<���<U��<���<J��<���<U��<���<e��<J��<���<b��<s��<R��<~��<���<`   `   ^��<���<���<���<���<O��<r��<4��<Y��<~��<N��<x��<A��<x��<N��<~��<Y��<4��<r��<O��<���<���<���<���<`   `   P��<b��<g��<���<Έ�<���<���<_��<c��<s��<j��<N��<��<N��<j��<s��<c��<_��<���<���<Έ�<���<g��<b��<`   `   ���<q��<���<���<���<���<r��<?��<[��<^��<R��<p��<T��<p��<R��<^��<[��<?��<r��<���<���<���<���<q��<`   `   ���<x��<���<Z��<c��<s��<C��<��<*��<s��<Z��<y��<��<y��<Z��<s��<*��<��<C��<s��<c��<Z��<���<x��<`   `   ���<t��<j��<g��<���<r��<w��<p��<��<a��<|��<i��<7��<i��<|��<a��<��<p��<w��<r��<���<g��<j��<t��<`   `   Ĉ�<|��<Y��<s��<���<Y��<���<���<.��<5��<]��<���<_��<���<]��<5��<.��<���<���<Y��<���<s��<Y��<|��<`   `   ���<V��<~��<q��<��<B��<X��<;��<]��<o��<D��<W��<n��<W��<D��<o��<]��<;��<X��<B��<��<q��<~��<V��<`   `   \��<-��<���<���<"��<���<���<`��<{��<���<W��<@��<u��<@��<W��<���<{��<`��<���<���<"��<���<���<-��<`   `   ���<S��<X��<���<g��<���<{��<���<���<c��<|��<���<Έ�<���<|��<c��<���<���<{��<���<g��<���<X��<S��<`   `   ���<���<O��<t��<e��<E��<8��<���<���<r��<���<���<b��<���<���<r��<���<���<8��<E��<e��<t��<O��<���<`   `   ~��<Z��<j��<���<n��<~��<���<���<���<���<���<���<:��<���<���<���<���<���<���<~��<n��<���<j��<Z��<`   `   W��<4��<z��<���<y��<u��<j��<f��<g��<\��<���<و�<���<و�<���<\��<g��<f��<j��<u��<y��<���<z��<4��<`   `   ���<c��<w��<���<���<���<R��<}��<���<c��<���<���<$��<���<���<c��<���<}��<R��<���<���<���<w��<c��<`   `   ���<���<f��<s��<���<w��<p��<���<���<���<���<���<��<���<���<���<���<���<p��<w��<���<s��<f��<���<`   `   ��<o��<W��<|��<���<E��<���<e��<`��<���<Ĉ�<Ɉ�<���<Ɉ�<Ĉ�<���<`��<e��<���<E��<���<|��<W��<o��<`   `   ��<���<���<c��<���<d��<È�<���<���<ƈ�<Y��<���<��<���<Y��<ƈ�<���<���<È�<d��<���<c��<���<���<`   `   G��<���<���<g��<���<���<��<W��<���<���<,��<x��<���<x��<,��<���<���<W��<��<���<���<g��<���<���<`   `   {��<&��<w��<���<���<���<E��<M��<���<ш�<���<���<H��<���<���<ш�<���<M��<E��<���<���<���<w��<&��<`   `   ˈ�<8��<q��<}��<���<���<���<���<���<���<؈�<���<���<���<؈�<���<���<���<���<���<���<}��<q��<8��<`   `   c��<��<{��<z��<j��<��<���<͈�<>��<2��<���<���<Q��<���<���<2��<>��<͈�<���<��<j��<z��<{��<��<`   `   -��<��<l��<���<���<���<Q��<���<y��<O��<���<���</��<���<���<O��<y��<���<Q��<���<���<���<l��<��<`   `   T��<y��<q��<Q��<W��<���<R��<���<��<���<͈�<���<���<���<͈�<���<��<���<R��<���<W��<Q��<q��<y��<`   `   ��<���<v��<b��<U��<���<���<���<���<h��<_��<j��<���<j��<_��<h��<���<���<���<���<U��<b��<v��<���<`   `   J��<���<U��<���<e��<J��<���<b��<s��<R��<~��<���<���<���<~��<R��<s��<b��<���<J��<e��<���<U��<���<`   `   A��<x��<N��<~��<Y��<4��<r��<O��<���<���<���<���<^��<���<���<���<���<O��<r��<4��<Y��<~��<N��<x��<`   `   ���<
��<��<��<��<7��<��<��<Ɇ�<ӆ�<��<��<1��<��<��<ӆ�<Ɇ�<��<��<7��<��<��<��<
��<`   `   ��<��<,��<��<+��<V��<���<(��<��<��<��<��<B��<��<��<��<��<(��<���<V��<+��<��<,��<��<`   `   І�<Ɇ�<��<��< ��<M��<���<4��<��<-��<5��<��<7��<��<5��<-��<��<4��<���<M��< ��<��<��<Ɇ�<`   `   4��<��<���<��<7��<7��<��<��<Ɔ�<���<��<��<��<��<��<���<Ɔ�<��<��<7��<7��<��<���<��<`   `   <��<��<	��<F��<G��<��<)��<C��<��<%��<%��<��<��<��<%��<%��<��<C��<)��<��<G��<F��<	��<��<`   `   ��<��<��<)��<��<��<��<9��<)��<E��<%��<��<��<��<%��<E��<)��<9��<��<��<��<)��<��<��<`   `   ��<'��<$��<���<��</��<���<��<M��<��<��<>��<��<>��<��<��<M��<��<���</��<��<���<$��<'��<`   `   φ�<��< ��<���<��<8��<��<��<\��< ��<	��<N��<��<N��<	��< ��<\��<��<��<8��<��<���< ��<��<`   `   ���<��<��<��<��<��<6��</��<'��<���<(��<��<���<��<(��<���<'��</��<6��<��<��<��<��<��<`   `   G��<��<��<+��<��<��<8��<5��<��<��<#��<��<	��<��<#��<��<��<5��<8��<��<��<+��<��<��<`   `   :��<��<��<3��<'��<��<��<��<��<��<��<:��<M��<:��<��<��<��<��<��<��<'��<3��<��<��<`   `   M��<,��<)��<!��<`��<G��<)��<F��<��<���<��<	��<ۆ�<	��<��<���<��<F��<)��<G��<`��<!��<)��<,��<`   `   v��<_��<<��<���<>��<&��<?��<M��<���<��<*��<<��<���<<��<*��<��<���<M��<?��<&��<>��<���<<��<_��<`   `   ��<��<+��<��<?��<,��<3��<��<��<:��<
��<<��<3��<<��<
��<:��<��<��<3��<,��<?��<��<+��<��<`   `   4��<+��<0��<6��<;��<>��<M��<��<��<.��<ņ�<���<��<���<ņ�<.��<��<��<M��<>��<;��<6��<0��<+��<`   `   Q��<���<J��<��<��<��<@��<��<��<��<��<!��<b��<!��<��<��<��<��<@��<��<��<��<J��<���<`   `   ӆ�<d��<2��<��<E��<5��<:��<���<Ն�<��<:��<��<<��<��<:��<��<Ն�<���<:��<5��<E��<��<2��<d��<`   `   9��<`��<��<C��<>��<��<0��<��<��<��< ��<��<��<��< ��<��<��<��<0��<��<>��<C��<��<`��<`   `   |��<@��<���<m��<+��<��<��<��<��<��<)��<8��<W��<8��<)��<��<��<��<��<��<+��<m��<���<@��<`   `   ��<��<:��<a��<3��<6��<"��<��<��<��<0��<3��<��<3��<0��<��<��<��<"��<6��<3��<a��<:��<��<`   `   E��<?��<V��<��<��<#��<��<���<!��<	��<��<��<��<��<��<	��<!��<���<��<#��<��<��<V��<?��<`   `   W��<��< ��<��<��<��<��<���<��<��<ֆ�<��<��<��<ֆ�<��<��<���<��<��<��<��< ��<��<`   `   G��<��<@��<F��<K��<(��<��< ��<��<I��<���<��<���<��<���<I��<��< ��<��<(��<K��<F��<@��<��<`   `   J��<@��<X��<��<��<��<$��<2��<��<'��<܆�<ц�<@��<ц�<܆�<'��<��<2��<$��<��<��<��<X��<@��<`   `   1��<��<��<ӆ�<Ɇ�<��<��<7��<��<��<��<
��<���<
��<��<��<��<7��<��<��<Ɇ�<ӆ�<��<��<`   `   B��<��<��<��<��<(��<���<V��<+��<��<,��<��<��<��<,��<��<+��<V��<���<(��<��<��<��<��<`   `   7��<��<5��<-��<��<4��<���<M��< ��<��<��<Ɇ�<І�<Ɇ�<��<��< ��<M��<���<4��<��<-��<5��<��<`   `   ��<��<��<���<Ɔ�<��<��<7��<7��<��<���<��<4��<��<���<��<7��<7��<��<��<Ɔ�<���<��<��<`   `   ��<��<%��<%��<��<C��<)��<��<G��<F��<	��<��<<��<��<	��<F��<G��<��<)��<C��<��<%��<%��<��<`   `   ��<��<%��<E��<)��<9��<��<��<��<)��<��<��<��<��<��<)��<��<��<��<9��<)��<E��<%��<��<`   `   ��<>��<��<��<M��<��<���</��<��<���<$��<'��<��<'��<$��<���<��</��<���<��<M��<��<��<>��<`   `   ��<N��<	��< ��<\��<��<��<8��<��<���< ��<��<φ�<��< ��<���<��<8��<��<��<\��< ��<	��<N��<`   `   ���<��<(��<���<'��</��<6��<��<��<��<��<��<���<��<��<��<��<��<6��</��<'��<���<(��<��<`   `   	��<��<#��<��<��<5��<8��<��<��<+��<��<��<G��<��<��<+��<��<��<8��<5��<��<��<#��<��<`   `   M��<:��<��<��<��<��<��<��<'��<3��<��<��<:��<��<��<3��<'��<��<��<��<��<��<��<:��<`   `   ۆ�<	��<��<���<��<F��<)��<G��<`��<!��<)��<,��<M��<,��<)��<!��<`��<G��<)��<F��<��<���<��<	��<`   `   ���<<��<*��<��<���<M��<?��<&��<>��<���<<��<_��<v��<_��<<��<���<>��<&��<?��<M��<���<��<*��<<��<`   `   3��<<��<
��<:��<��<��<3��<,��<?��<��<+��<��<��<��<+��<��<?��<,��<3��<��<��<:��<
��<<��<`   `   ��<���<ņ�<.��<��<��<M��<>��<;��<6��<0��<+��<4��<+��<0��<6��<;��<>��<M��<��<��<.��<ņ�<���<`   `   b��<!��<��<��<��<��<@��<��<��<��<J��<���<Q��<���<J��<��<��<��<@��<��<��<��<��<!��<`   `   <��<��<:��<��<Ն�<���<:��<5��<E��<��<2��<d��<ӆ�<d��<2��<��<E��<5��<:��<���<Ն�<��<:��<��<`   `   ��<��< ��<��<��<��<0��<��<>��<C��<��<`��<9��<`��<��<C��<>��<��<0��<��<��<��< ��<��<`   `   W��<8��<)��<��<��<��<��<��<+��<m��<���<@��<|��<@��<���<m��<+��<��<��<��<��<��<)��<8��<`   `   ��<3��<0��<��<��<��<"��<6��<3��<a��<:��<��<��<��<:��<a��<3��<6��<"��<��<��<��<0��<3��<`   `   ��<��<��<	��<!��<���<��<#��<��<��<V��<?��<E��<?��<V��<��<��<#��<��<���<!��<	��<��<��<`   `   ��<��<ֆ�<��<��<���<��<��<��<��< ��<��<W��<��< ��<��<��<��<��<���<��<��<ֆ�<��<`   `   ���<��<���<I��<��< ��<��<(��<K��<F��<@��<��<G��<��<@��<F��<K��<(��<��< ��<��<I��<���<��<`   `   @��<ц�<܆�<'��<��<2��<$��<��<��<��<X��<@��<J��<@��<X��<��<��<��<$��<2��<��<'��<܆�<ц�<`   `   ���<���<Ѕ�<���<���<���<���<���<��<��<��<��<߅�<��<��<��<��<���<���<���<���<���<Ѕ�<���<`   `   ���<���<؅�<Å�<���<���<���<���<���<��<ʅ�<߅�<���<߅�<ʅ�<��<���<���<���<���<���<Å�<؅�<���<`   `   ��<Ѕ�<��<���<���<���<��<΅�<م�<݅�<���<Ӆ�<���<Ӆ�<���<݅�<م�<΅�<��<���<���<���<��<Ѕ�<`   `   ��<Ʌ�<˅�<���<���<���<���<Ʌ�<Յ�<��<υ�<��<Ѕ�<��<υ�<��<Յ�<Ʌ�<���<���<���<���<˅�<Ʌ�<`   `   ���<���<ą�<���<���<���<���<ǅ�<���<Ѕ�<х�<܅�<���<܅�<х�<Ѕ�<���<ǅ�<���<���<���<���<ą�<���<`   `   ���<Ʌ�<ƅ�<���<���<��<؅�<̅�<Յ�<���<���<ׅ�<���<ׅ�<���<���<Յ�<̅�<؅�<��<���<���<ƅ�<Ʌ�<`   `   ���<���<���<���<���<҅�<���<���<݅�<���<���<��<���<��<���<���<݅�<���<���<҅�<���<���<���<���<`   `   ʅ�<ƅ�<���<���<ą�<���<߅�<Ņ�<���<���<ۅ�<��<���<��<ۅ�<���<���<Ņ�<߅�<���<ą�<���<���<ƅ�<`   `   ��<��<���<���<��<҅�<��<Ѕ�<���<څ�<��<���<΅�<���<��<څ�<���<Ѕ�<��<҅�<��<���<���<��<`   `   ��<օ�<���<Ӆ�<���<���<���<���<Ѕ�<Յ�<���<���<ׅ�<���<���<Յ�<Ѕ�<���<���<���<���<Ӆ�<���<օ�<`   `   ���<���<��<��<ą�<��<Յ�<���<��<Ʌ�<���<��<օ�<��<���<Ʌ�<��<���<Յ�<��<ą�<��<��<���<`   `   ���<���<���<���<���<���<ޅ�<���<˅�<��<�<Ӆ�<���<Ӆ�<�<��<˅�<���<ޅ�<���<���<���<���<���<`   `   *��<���<ʅ�<��<���<���<���<΅�<���<��<���<���<���<���<���<��<���<΅�<���<���<���<��<ʅ�<���<`   `   ��<���<��<Ӆ�< ��<Ӆ�<���<��<���<΅�<х�<΅�<߅�<΅�<х�<΅�<���<��<���<Ӆ�< ��<Ӆ�<��<���<`   `   ���<���<��<˅�<΅�<���<���<	��<Յ�<��<��<���<���<���<��<��<Յ�<	��<���<���<΅�<˅�<��<���<`   `   օ�<х�<��<��<ۅ�<߅�<���<��<���<م�<ą�<���<���<���<ą�<م�<���<��<���<߅�<ۅ�<��<��<х�<`   `   ��<օ�<څ�<΅�<ۅ�<��<���<݅�<��<���<���<څ�<���<څ�<���<���<��<݅�<���<��<ۅ�<΅�<څ�<օ�<`   `   ǅ�<���<���<���<���<���<�<ƅ�<��<΅�<̅�<ʅ�<n��<ʅ�<̅�<΅�<��<ƅ�<�<���<���<���<���<���<`   `   ��<߅�<ׅ�<%��<��<���<���<�<���<���<���<�<���<�<���<���<���<�<���<���<��<%��<ׅ�<߅�<`   `   ��<��<���<��<��<ޅ�<��<���<���<���<���<���<���<���<���<���<���<���<��<ޅ�<��<��<���<��<`   `   օ�<ą�<���<���<���<��<#��<Յ�<څ�<���<���<���<���<���<���<���<څ�<Յ�<#��<��<���<���<���<ą�<`   `   ��<���<��<��<ͅ�<΅�<օ�<܅�<ƅ�<���<���<΅�<��<΅�<���<���<ƅ�<܅�<օ�<΅�<ͅ�<��<��<���<`   `   ��<���<΅�<؅�<���<ƅ�<���<��<���<���<��<ͅ�<���<ͅ�<��<���<���<��<���<ƅ�<���<؅�<΅�<���<`   `   ͅ�<���<���<Ʌ�<ׅ�<
��<���<��<���<���<��<���<���<���<��<���<���<��<���<
��<ׅ�<Ʌ�<���<���<`   `   ߅�<��<��<��<��<���<���<���<���<���<Ѕ�<���<���<���<Ѕ�<���<���<���<���<���<��<��<��<��<`   `   ���<߅�<ʅ�<��<���<���<���<���<���<Å�<؅�<���<���<���<؅�<Å�<���<���<���<���<���<��<ʅ�<߅�<`   `   ���<Ӆ�<���<݅�<م�<΅�<��<���<���<���<��<Ѕ�<��<Ѕ�<��<���<���<���<��<΅�<م�<݅�<���<Ӆ�<`   `   Ѕ�<��<υ�<��<Յ�<Ʌ�<���<���<���<���<˅�<Ʌ�<��<Ʌ�<˅�<���<���<���<���<Ʌ�<Յ�<��<υ�<��<`   `   ���<܅�<х�<Ѕ�<���<ǅ�<���<���<���<���<ą�<���<���<���<ą�<���<���<���<���<ǅ�<���<Ѕ�<х�<܅�<`   `   ���<ׅ�<���<���<Յ�<̅�<؅�<��<���<���<ƅ�<Ʌ�<���<Ʌ�<ƅ�<���<���<��<؅�<̅�<Յ�<���<���<ׅ�<`   `   ���<��<���<���<݅�<���<���<҅�<���<���<���<���<���<���<���<���<���<҅�<���<���<݅�<���<���<��<`   `   ���<��<ۅ�<���<���<Ņ�<߅�<���<ą�<���<���<ƅ�<ʅ�<ƅ�<���<���<ą�<���<߅�<Ņ�<���<���<ۅ�<��<`   `   ΅�<���<��<څ�<���<Ѕ�<��<҅�<��<���<���<��<��<��<���<���<��<҅�<��<Ѕ�<���<څ�<��<���<`   `   ׅ�<���<���<Յ�<Ѕ�<���<���<���<���<Ӆ�<���<օ�<��<օ�<���<Ӆ�<���<���<���<���<Ѕ�<Յ�<���<���<`   `   օ�<��<���<Ʌ�<��<���<Յ�<��<ą�<��<��<���<���<���<��<��<ą�<��<Յ�<���<��<Ʌ�<���<��<`   `   ���<Ӆ�<�<��<˅�<���<ޅ�<���<���<���<���<���<���<���<���<���<���<���<ޅ�<���<˅�<��<�<Ӆ�<`   `   ���<���<���<��<���<΅�<���<���<���<��<ʅ�<���<*��<���<ʅ�<��<���<���<���<΅�<���<��<���<���<`   `   ߅�<΅�<х�<΅�<���<��<���<Ӆ�< ��<Ӆ�<��<���<��<���<��<Ӆ�< ��<Ӆ�<���<��<���<΅�<х�<΅�<`   `   ���<���<��<��<Յ�<	��<���<���<΅�<˅�<��<���<���<���<��<˅�<΅�<���<���<	��<Յ�<��<��<���<`   `   ���<���<ą�<م�<���<��<���<߅�<ۅ�<��<��<х�<օ�<х�<��<��<ۅ�<߅�<���<��<���<م�<ą�<���<`   `   ���<څ�<���<���<��<݅�<���<��<ۅ�<΅�<څ�<օ�<��<օ�<څ�<΅�<ۅ�<��<���<݅�<��<���<���<څ�<`   `   n��<ʅ�<̅�<΅�<��<ƅ�<�<���<���<���<���<���<ǅ�<���<���<���<���<���<�<ƅ�<��<΅�<̅�<ʅ�<`   `   ���<�<���<���<���<�<���<���<��<%��<ׅ�<߅�<��<߅�<ׅ�<%��<��<���<���<�<���<���<���<�<`   `   ���<���<���<���<���<���<��<ޅ�<��<��<���<��<��<��<���<��<��<ޅ�<��<���<���<���<���<���<`   `   ���<���<���<���<څ�<Յ�<#��<��<���<���<���<ą�<օ�<ą�<���<���<���<��<#��<Յ�<څ�<���<���<���<`   `   ��<΅�<���<���<ƅ�<܅�<օ�<΅�<ͅ�<��<��<���<��<���<��<��<ͅ�<΅�<օ�<܅�<ƅ�<���<���<΅�<`   `   ���<ͅ�<��<���<���<��<���<ƅ�<���<؅�<΅�<���<��<���<΅�<؅�<���<ƅ�<���<��<���<���<��<ͅ�<`   `   ���<���<��<���<���<��<���<
��<ׅ�<Ʌ�<���<���<ͅ�<���<���<Ʌ�<ׅ�<
��<���<��<���<���<��<���<`   `   s��<���<_��<{��<���<��<���<���<���<���<t��<���<x��<���<t��<���<���<���<���<��<���<{��<_��<���<`   `   ���<���<S��<���<���<a��<���<V��<h��<\��<U��<���<Z��<���<U��<\��<h��<V��<���<a��<���<���<S��<���<`   `   n��<x��<^��<���<���<d��<���<T��<��<m��<b��<Ą�<c��<Ą�<b��<m��<��<T��<���<d��<���<���<^��<x��<`   `   X��<e��<���<���<���<���<���<���<���<���<e��<���<x��<���<e��<���<���<���<���<���<���<���<���<e��<`   `   ���<���<���<x��<u��<���<���<w��<���<���<Y��<z��<���<z��<Y��<���<���<w��<���<���<u��<x��<���<���<`   `   ���<~��<���<���<���<���<���<a��<p��<���<���<���<���<���<���<���<p��<a��<���<���<���<���<���<~��<`   `   y��<X��<f��<Ä�<���<a��<���<���<}��<˄�<���<j��<���<j��<���<˄�<}��<���<���<a��<���<Ä�<f��<X��<`   `   t��<y��<r��<���<y��<`��<���<���<m��<���<x��<1��<���<1��<x��<���<m��<���<���<`��<y��<���<r��<y��<`   `   E��<���<���<V��<���<���<h��<���<j��<���<d��<m��<#��<m��<d��<���<j��<���<h��<���<���<V��<���<���<`   `   +��<���<���<S��<���<u��<5��<���<���<���<���<k��<���<k��<���<���<���<���<5��<u��<���<S��<���<���<`   `   ���<҄�<���<\��<���<u��<���<Ʉ�<���<e��<���<k��<��<k��<���<e��<���<Ʉ�<���<u��<���<\��<���<҄�<`   `   ���<���<���<}��<���<���<���<i��<���<���<���<ń�<���<ń�<���<���<���<i��<���<���<���<}��<���<���<`   `   1��<j��<���<���<���<���<���<f��<���<���<[��<���<Ä�<���<[��<���<���<f��<���<���<���<���<���<j��<`   `   ؄�<҄�<Ǆ�<���<���<Є�<���<���<|��<`��<w��<p��<z��<p��<w��<`��<|��<���<���<Є�<���<���<Ǆ�<҄�<`   `   ��<���<���<_��<w��<���<���<z��<2��<_��<���<���<{��<���<���<_��<2��<z��<���<���<w��<_��<���<���<`   `   ���<#��<;��<���<���<���<y��<t��<~��<���<}��<���<i��<���<}��<���<~��<t��<y��<���<���<���<;��<#��<`   `   !��<���<���<ل�<���<b��<n��<m��<~��<|��<Y��<���<���<���<Y��<|��<~��<m��<n��<b��<���<ل�<���<���<`   `   ���<���<��<���<���<���<���<i��<[��<���<���<���<���<���<���<���<[��<i��<���<���<���<���<��<���<`   `   ��<���<��<7��<���<��<���<���<s��<���<���<z��<���<z��<���<���<s��<���<���<��<���<7��<��<���<`   `   q��<Ä�<���<Z��<���<Z��<O��<���<d��<{��<���<���<���<���<���<{��<d��<���<O��<Z��<���<Z��<���<Ä�<`   `   W��<���<���<���<҄�<T��<?��<q��<c��<z��<���<���<}��<���<���<z��<c��<q��<?��<T��<҄�<���<���<���<`   `   h��<���<���<���<Ǆ�<���<���<v��<���<���<���<^��<l��<^��<���<���<���<v��<���<���<Ǆ�<���<���<���<`   `   ���<Є�<���<Q��<X��<���<���<r��<���<y��<n��<l��<���<l��<n��<y��<���<r��<���<���<X��<Q��<���<Є�<`   `   ���<���<���<���<i��<n��<o��<p��<���<w��<y��<���<���<���<y��<w��<���<p��<o��<n��<i��<���<���<���<`   `   x��<���<t��<���<���<���<���<��<���<{��<_��<���<s��<���<_��<{��<���<��<���<���<���<���<t��<���<`   `   Z��<���<U��<\��<h��<V��<���<a��<���<���<S��<���<���<���<S��<���<���<a��<���<V��<h��<\��<U��<���<`   `   c��<Ą�<b��<m��<��<T��<���<d��<���<���<^��<x��<n��<x��<^��<���<���<d��<���<T��<��<m��<b��<Ą�<`   `   x��<���<e��<���<���<���<���<���<���<���<���<e��<X��<e��<���<���<���<���<���<���<���<���<e��<���<`   `   ���<z��<Y��<���<���<w��<���<���<u��<x��<���<���<���<���<���<x��<u��<���<���<w��<���<���<Y��<z��<`   `   ���<���<���<���<p��<a��<���<���<���<���<���<~��<���<~��<���<���<���<���<���<a��<p��<���<���<���<`   `   ���<j��<���<˄�<}��<���<���<a��<���<Ä�<f��<X��<y��<X��<f��<Ä�<���<a��<���<���<}��<˄�<���<j��<`   `   ���<1��<x��<���<m��<���<���<`��<y��<���<r��<y��<t��<y��<r��<���<y��<`��<���<���<m��<���<x��<1��<`   `   #��<m��<d��<���<j��<���<h��<���<���<V��<���<���<E��<���<���<V��<���<���<h��<���<j��<���<d��<m��<`   `   ���<k��<���<���<���<���<5��<u��<���<S��<���<���<+��<���<���<S��<���<u��<5��<���<���<���<���<k��<`   `   ��<k��<���<e��<���<Ʉ�<���<u��<���<\��<���<҄�<���<҄�<���<\��<���<u��<���<Ʉ�<���<e��<���<k��<`   `   ���<ń�<���<���<���<i��<���<���<���<}��<���<���<���<���<���<}��<���<���<���<i��<���<���<���<ń�<`   `   Ä�<���<[��<���<���<f��<���<���<���<���<���<j��<1��<j��<���<���<���<���<���<f��<���<���<[��<���<`   `   z��<p��<w��<`��<|��<���<���<Є�<���<���<Ǆ�<҄�<؄�<҄�<Ǆ�<���<���<Є�<���<���<|��<`��<w��<p��<`   `   {��<���<���<_��<2��<z��<���<���<w��<_��<���<���<��<���<���<_��<w��<���<���<z��<2��<_��<���<���<`   `   i��<���<}��<���<~��<t��<y��<���<���<���<;��<#��<���<#��<;��<���<���<���<y��<t��<~��<���<}��<���<`   `   ���<���<Y��<|��<~��<m��<n��<b��<���<ل�<���<���<!��<���<���<ل�<���<b��<n��<m��<~��<|��<Y��<���<`   `   ���<���<���<���<[��<i��<���<���<���<���<��<���<���<���<��<���<���<���<���<i��<[��<���<���<���<`   `   ���<z��<���<���<s��<���<���<��<���<7��<��<���<��<���<��<7��<���<��<���<���<s��<���<���<z��<`   `   ���<���<���<{��<d��<���<O��<Z��<���<Z��<���<Ä�<q��<Ä�<���<Z��<���<Z��<O��<���<d��<{��<���<���<`   `   }��<���<���<z��<c��<q��<?��<T��<҄�<���<���<���<W��<���<���<���<҄�<T��<?��<q��<c��<z��<���<���<`   `   l��<^��<���<���<���<v��<���<���<Ǆ�<���<���<���<h��<���<���<���<Ǆ�<���<���<v��<���<���<���<^��<`   `   ���<l��<n��<y��<���<r��<���<���<X��<Q��<���<Є�<���<Є�<���<Q��<X��<���<���<r��<���<y��<n��<l��<`   `   ���<���<y��<w��<���<p��<o��<n��<i��<���<���<���<���<���<���<���<i��<n��<o��<p��<���<w��<y��<���<`   `   ��<W��<X��<B��<��<R��<X��<,��<@��< ��<7��<J��<[��<J��<7��< ��<@��<,��<X��<R��<��<B��<X��<W��<`   `   5��<t��<_��<I��<E��<d��<L��<h��<���<t��<z��<Z��<_��<Z��<z��<t��<���<h��<L��<d��<E��<I��<_��<t��<`   `   -��<^��<O��<N��<T��<=��<��<F��<t��<���<���<L��<Q��<L��<���<���<t��<F��<��<=��<T��<N��<O��<^��<`   `   8��<D��<>��<M��<[��<G��<4��<G��<��<A��<p��<2��<:��<2��<p��<A��<��<G��<4��<G��<[��<M��<>��<D��<`   `   ���<U��<5��<J��<D��<4��</��<e��<Q��<\��<z��<H��<L��<H��<z��<\��<Q��<e��</��<4��<D��<J��<5��<U��<`   `   L��<9��<:��<N��<5��<.��<:��<x��<h��<C��<C��<<��<c��<<��<C��<C��<h��<x��<:��<.��<5��<N��<:��<9��<`   `   A��<f��<c��<>��<D��<U��<F��<c��<=��<��<B��<Z��<���<Z��<B��<��<=��<c��<F��<U��<D��<>��<c��<f��<`   `   }��<���<h��<+��<V��<���<,��<A��<N��<(��<]��<W��<L��<W��<]��<(��<N��<A��<,��<���<V��<+��<h��<���<`   `   ��<V��<_��<Y��<E��<���<_��<a��<s��<1��<c��<P��<��<P��<c��<1��<s��<a��<_��<���<E��<Y��<_��<V��<`   `   u��<6��<S��<���<S��<T��<���<c��<A��<E��<���<���<I��<���<���<E��<A��<c��<���<T��<S��<���<S��<6��<`   `   W��<=��<��<���<���<,��<_��<U��<*��<S��<c��<V��<Y��<V��<c��<S��<*��<U��<_��<,��<���<���<��<=��<`   `   c��<���<)��<R��<���<8��<M��<U��<F��<>��<B��<3��<G��<3��<B��<>��<F��<U��<M��<8��<���<R��<)��<���<`   `   C��<���<J��<T��<<��<4��<T��<M��<a��<<��<r��<@��<"��<@��<r��<<��<a��<M��<T��<4��<<��<T��<J��<���<`   `   ��<@��</��<x��<%��<��<<��<J��<���<e��<x��<F��<>��<F��<x��<e��<���<J��<<��<��<%��<x��</��<@��<`   `   ��<o��<t��<���<i��<C��<d��<H��<���<l��<4��<M��<���<M��<4��<l��<���<H��<d��<C��<i��<���<t��<o��<`   `   (��<���<���<Z��<Z��<n��<���<\��<f��<x��</��<I��<e��<I��</��<x��<f��<\��<���<n��<Z��<Z��<���<���<`   `   D��<`��<`��<��<=��<)��<���<���<Y��<~��<O��<J��<��<J��<O��<~��<Y��<���<���<)��<=��<��<`��<`��<`   `   ���<)��<(��<I��<���<'��<A��<���<+��<X��<4��<3��<-��<3��<4��<X��<+��<���<A��<'��<���<I��<(��<)��<`   `   ���<4��<-��<Q��<y��<=��<$��<h��<0��<h��<G��<:��<a��<:��<G��<h��<0��<h��<$��<=��<y��<Q��<-��<4��<`   `   ���<M��<X��<��<^��<o��<_��<���<y��<O��<Q��<O��<f��<O��<Q��<O��<y��<���<_��<o��<^��<��<X��<M��<`   `   ���<f��<I��<v��<D��<n��<z��<~��<u��<��<E��<S��<J��<S��<E��<��<u��<~��<z��<n��<D��<v��<I��<f��<`   `   C��<c��<��<'��<��<7��<g��<B��<c��<J��<W��<M��<Z��<M��<W��<J��<c��<B��<g��<7��<��<'��<��<c��<`   `   ���<S��<b��<���<���<b��<���<G��<\��<v��<:��<:��<{��<:��<:��<v��<\��<G��<���<b��<���<���<b��<S��<`   `   3��<Y��<y��<���<}��<;��<g��<3��<��<P��<4��<D��<^��<D��<4��<P��<��<3��<g��<;��<}��<���<y��<Y��<`   `   [��<J��<7��< ��<@��<,��<X��<R��<��<B��<X��<W��<��<W��<X��<B��<��<R��<X��<,��<@��< ��<7��<J��<`   `   _��<Z��<z��<t��<���<h��<L��<d��<E��<I��<_��<t��<5��<t��<_��<I��<E��<d��<L��<h��<���<t��<z��<Z��<`   `   Q��<L��<���<���<t��<F��<��<=��<T��<N��<O��<^��<-��<^��<O��<N��<T��<=��<��<F��<t��<���<���<L��<`   `   :��<2��<p��<A��<��<G��<4��<G��<[��<M��<>��<D��<8��<D��<>��<M��<[��<G��<4��<G��<��<A��<p��<2��<`   `   L��<H��<z��<\��<Q��<e��</��<4��<D��<J��<5��<U��<���<U��<5��<J��<D��<4��</��<e��<Q��<\��<z��<H��<`   `   c��<<��<C��<C��<h��<x��<:��<.��<5��<N��<:��<9��<L��<9��<:��<N��<5��<.��<:��<x��<h��<C��<C��<<��<`   `   ���<Z��<B��<��<=��<c��<F��<U��<D��<>��<c��<f��<A��<f��<c��<>��<D��<U��<F��<c��<=��<��<B��<Z��<`   `   L��<W��<]��<(��<N��<A��<,��<���<V��<+��<h��<���<}��<���<h��<+��<V��<���<,��<A��<N��<(��<]��<W��<`   `   ��<P��<c��<1��<s��<a��<_��<���<E��<Y��<_��<V��<��<V��<_��<Y��<E��<���<_��<a��<s��<1��<c��<P��<`   `   I��<���<���<E��<A��<c��<���<T��<S��<���<S��<6��<u��<6��<S��<���<S��<T��<���<c��<A��<E��<���<���<`   `   Y��<V��<c��<S��<*��<U��<_��<,��<���<���<��<=��<W��<=��<��<���<���<,��<_��<U��<*��<S��<c��<V��<`   `   G��<3��<B��<>��<F��<U��<M��<8��<���<R��<)��<���<c��<���<)��<R��<���<8��<M��<U��<F��<>��<B��<3��<`   `   "��<@��<r��<<��<a��<M��<T��<4��<<��<T��<J��<���<C��<���<J��<T��<<��<4��<T��<M��<a��<<��<r��<@��<`   `   >��<F��<x��<e��<���<J��<<��<��<%��<x��</��<@��<��<@��</��<x��<%��<��<<��<J��<���<e��<x��<F��<`   `   ���<M��<4��<l��<���<H��<d��<C��<i��<���<t��<o��<��<o��<t��<���<i��<C��<d��<H��<���<l��<4��<M��<`   `   e��<I��</��<x��<f��<\��<���<n��<Z��<Z��<���<���<(��<���<���<Z��<Z��<n��<���<\��<f��<x��</��<I��<`   `   ��<J��<O��<~��<Y��<���<���<)��<=��<��<`��<`��<D��<`��<`��<��<=��<)��<���<���<Y��<~��<O��<J��<`   `   -��<3��<4��<X��<+��<���<A��<'��<���<I��<(��<)��<���<)��<(��<I��<���<'��<A��<���<+��<X��<4��<3��<`   `   a��<:��<G��<h��<0��<h��<$��<=��<y��<Q��<-��<4��<���<4��<-��<Q��<y��<=��<$��<h��<0��<h��<G��<:��<`   `   f��<O��<Q��<O��<y��<���<_��<o��<^��<��<X��<M��<���<M��<X��<��<^��<o��<_��<���<y��<O��<Q��<O��<`   `   J��<S��<E��<��<u��<~��<z��<n��<D��<v��<I��<f��<���<f��<I��<v��<D��<n��<z��<~��<u��<��<E��<S��<`   `   Z��<M��<W��<J��<c��<B��<g��<7��<��<'��<��<c��<C��<c��<��<'��<��<7��<g��<B��<c��<J��<W��<M��<`   `   {��<:��<:��<v��<\��<G��<���<b��<���<���<b��<S��<���<S��<b��<���<���<b��<���<G��<\��<v��<:��<:��<`   `   ^��<D��<4��<P��<��<3��<g��<;��<}��<���<y��<Y��<3��<Y��<y��<���<}��<;��<g��<3��<��<P��<4��<D��<`   `   ��<��<.��<U��<(��<@��<���<B��<��< ��<\��<��<^��<��<\��< ��<��<B��<���<@��<(��<U��<.��<��<`   `   "��<���<��<8��<��<S��<��<N��<$��<��<Z��<��<V��<��<Z��<��<$��<N��<��<S��<��<8��<��<���<`   `   K��<1��<+��<&��< ��<K��<(��<K��<���<��<��<��<���<��<��<��<���<K��<(��<K��< ��<&��<+��<1��<`   `   +��<?��<;��<��<	��<>��<J��<^��<#��<��<��<��<���<��<��<��<#��<^��<J��<>��<	��<��<;��<?��<`   `   ��<��<%��<>��<=��<=��<(��< ��<8��<5��<T��<X��<X��<X��<T��<5��<8��< ��<(��<=��<=��<>��<%��<��<`   `   ��<(��<+��<:��<;��<N��<A��<
��<-��<��<!��<��<��<��<!��<��<-��<
��<A��<N��<;��<:��<+��<(��<`   `   ��<J��<9��<��<"��<I��<T��<��<8��<7��<'��<!��<��<!��<'��<7��<8��<��<T��<I��<"��<��<9��<J��<`   `   ��<��<��<C��<K��<��<��<��<N��<:��<U��<h��<!��<h��<U��<:��<N��<��<��<��<K��<C��<��<��<`   `   /��<��<��<X��<��<���<��<��<a��<��<��<5��<���<5��<��<��<a��<��<��<���<��<X��<��<��<`   `   ���<M��<8��<*��<��<6��<T��<��<.��<,��<��<+��<(��<+��<��<,��<.��<��<T��<6��<��<*��<8��<M��<`   `   ��<��<K��<��<��<K��<#��<��<J��<y��<��<��<���<��<��<y��<J��<��<#��<K��<��<��<K��<��<`   `   ׁ�<��<]��<*��<��<-��<��<U��<h��<V��<.��<	��<K��<	��<.��<V��<h��<U��<��<-��<��<*��<]��<��<`   `   m��<g��<S��<T��<��<v��<a��<9��<���<��<`��<:��<A��<:��<`��<��<���<9��<a��<v��<��<T��<S��<g��<`   `   _��<A��<��<Z��<S��<l��<R��<
��<��<��<D��<$��<I��<$��<D��<��<��<
��<R��<l��<S��<Z��<��<A��<`   `   -��<T��<��<2��<O��<��< ��<1��<I��<��<��<��<-��<��<��<��<I��<1��< ��<��<O��<2��<��<T��<`   `   ��<z��<0��<��<@��<%��<��<���<��<���<F��<;��<��<;��<F��<���<��<���<��<%��<@��<��<0��<z��<`   `   ��<*��<>��<��<U��<d��<��<���< ��<��<V��<[��<��<[��<V��<��< ��<���<��<d��<U��<��<>��<*��<`   `   N��<7��<c��<e��<S��<N��<@��<N��<W��<)��<��<G��<6��<G��<��<)��<W��<N��<@��<N��<S��<e��<c��<7��<`   `   ���<J��<i��<b��<���<��<$��<��<��<(��<+��<A��<2��<A��<+��<(��<��<��<$��<��<���<b��<i��<J��<`   `   ���<��</��<=��<���<`��<<��<ԁ�<"��<>��<2��<��<���<��<2��<>��<"��<ԁ�<<��<`��<���<=��</��<��<`   `   ��<'��<G��<I��<��<z��<>��<��<<��<+��<(��<��<��<��<(��<+��<<��<��<>��<z��<��<I��<G��<'��<`   `   W��<h��<T��<Q��<��<��<��<��<��<��<P��<5��<'��<5��<P��<��<��<��<��<��<��<Q��<T��<h��<`   `   >��<,��<��<(��<E��<��<��<I��<��<��<<��<!��<��<!��<<��<��<��<I��<��<��<E��<(��<��<,��<`   `   w��<0��<��<��<!��<=��<��<O��<1��<6��<9��<2��<��<2��<9��<6��<1��<O��<��<=��<!��<��<��<0��<`   `   ^��<��<\��< ��<��<B��<���<@��<(��<U��<.��<��<��<��<.��<U��<(��<@��<���<B��<��< ��<\��<��<`   `   V��<��<Z��<��<$��<N��<��<S��<��<8��<��<���<"��<���<��<8��<��<S��<��<N��<$��<��<Z��<��<`   `   ���<��<��<��<���<K��<(��<K��< ��<&��<+��<1��<K��<1��<+��<&��< ��<K��<(��<K��<���<��<��<��<`   `   ���<��<��<��<#��<^��<J��<>��<	��<��<;��<?��<+��<?��<;��<��<	��<>��<J��<^��<#��<��<��<��<`   `   X��<X��<T��<5��<8��< ��<(��<=��<=��<>��<%��<��<��<��<%��<>��<=��<=��<(��< ��<8��<5��<T��<X��<`   `   ��<��<!��<��<-��<
��<A��<N��<;��<:��<+��<(��<��<(��<+��<:��<;��<N��<A��<
��<-��<��<!��<��<`   `   ��<!��<'��<7��<8��<��<T��<I��<"��<��<9��<J��<��<J��<9��<��<"��<I��<T��<��<8��<7��<'��<!��<`   `   !��<h��<U��<:��<N��<��<��<��<K��<C��<��<��<��<��<��<C��<K��<��<��<��<N��<:��<U��<h��<`   `   ���<5��<��<��<a��<��<��<���<��<X��<��<��</��<��<��<X��<��<���<��<��<a��<��<��<5��<`   `   (��<+��<��<,��<.��<��<T��<6��<��<*��<8��<M��<���<M��<8��<*��<��<6��<T��<��<.��<,��<��<+��<`   `   ���<��<��<y��<J��<��<#��<K��<��<��<K��<��<��<��<K��<��<��<K��<#��<��<J��<y��<��<��<`   `   K��<	��<.��<V��<h��<U��<��<-��<��<*��<]��<��<ׁ�<��<]��<*��<��<-��<��<U��<h��<V��<.��<	��<`   `   A��<:��<`��<��<���<9��<a��<v��<��<T��<S��<g��<m��<g��<S��<T��<��<v��<a��<9��<���<��<`��<:��<`   `   I��<$��<D��<��<��<
��<R��<l��<S��<Z��<��<A��<_��<A��<��<Z��<S��<l��<R��<
��<��<��<D��<$��<`   `   -��<��<��<��<I��<1��< ��<��<O��<2��<��<T��<-��<T��<��<2��<O��<��< ��<1��<I��<��<��<��<`   `   ��<;��<F��<���<��<���<��<%��<@��<��<0��<z��<��<z��<0��<��<@��<%��<��<���<��<���<F��<;��<`   `   ��<[��<V��<��< ��<���<��<d��<U��<��<>��<*��<��<*��<>��<��<U��<d��<��<���< ��<��<V��<[��<`   `   6��<G��<��<)��<W��<N��<@��<N��<S��<e��<c��<7��<N��<7��<c��<e��<S��<N��<@��<N��<W��<)��<��<G��<`   `   2��<A��<+��<(��<��<��<$��<��<���<b��<i��<J��<���<J��<i��<b��<���<��<$��<��<��<(��<+��<A��<`   `   ���<��<2��<>��<"��<ԁ�<<��<`��<���<=��</��<��<���<��</��<=��<���<`��<<��<ԁ�<"��<>��<2��<��<`   `   ��<��<(��<+��<<��<��<>��<z��<��<I��<G��<'��<��<'��<G��<I��<��<z��<>��<��<<��<+��<(��<��<`   `   '��<5��<P��<��<��<��<��<��<��<Q��<T��<h��<W��<h��<T��<Q��<��<��<��<��<��<��<P��<5��<`   `   ��<!��<<��<��<��<I��<��<��<E��<(��<��<,��<>��<,��<��<(��<E��<��<��<I��<��<��<<��<!��<`   `   ��<2��<9��<6��<1��<O��<��<=��<!��<��<��<0��<w��<0��<��<��<!��<=��<��<O��<1��<6��<9��<2��<`   `   7��<5��<��<��<��<��<��<(��<B��<a��<B��<��<���<��<B��<a��<B��<(��<��<��<��<��<��<5��<`   `   ;��<��<���<��<��<��<��<���<���<��<��<��<��<��<��<��<���<���<��<��<��<��<���<��<`   `   ��<���<��<=��<#��<��< ��<��<	��<)��<J��<=��<+��<=��<J��<)��<	��<��< ��<��<#��<=��<��<���<`   `   ���<���<���<��<��<���<��<���<T��<`��<(��<���<���<���<(��<`��<T��<���<��<���<��<��<���<���<`   `   ��<&��<��<���<��<���<��<��<��<��<ۀ�<��<Հ�<��<ۀ�<��<��<��<��<���<��<���<��<&��<`   `   4��<��<��<"��<��<��<	��<���<��<��<��<F��<$��<F��<��<��<��<���<	��<��<��<"��<��<��<`   `   1��<��<��<��<���<р�<��<��<��<I��<��<���<&��<���<��<I��<��<��<��<р�<���<��<��<��<`   `   ;��<D��<��<��<��<���<O��<$��<̀�<��<р�<��<I��<��<р�<��<̀�<$��<O��<���<��<��<��<D��<`   `   ��<3��<)��<��<@��<��<-��<+��<��<��<��<)��<K��<)��<��<��<��<+��<-��<��<@��<��<)��<3��<`   `   ���<��<��<݀�<F��<��<��<4��<��< ��<-��<2��<��<2��<-��< ��<��<4��<��<��<F��<݀�<��<��<`   `   ,��<-��<>��<���<M��<@��<��<A��<܀�<���<)��<��<Ԁ�<��<)��<���<܀�<A��<��<@��<M��<���<>��<-��<`   `   ]��<���<
��<��<"��<��<��</��<��<��<2��<��<��<��<2��<��<��</��<��<��<"��<��<
��<���<`   `   	��<ƀ�<���<��<���<��<̀�<��<7��<!��<���<���<&��<���<���<!��<7��<��<̀�<��<���<��<���<ƀ�<`   `   ��<*��<W��<��<��<��<���<���<5��<?��<���<��</��<��<���<?��<5��<���<���<��<��<��<W��<*��<`   `   ���<'��<2��<��<��<��<5��<<��<��<%��<J��<��<��<��<J��<%��<��<<��<5��<��<��<��<2��<'��<`   `   ?��<��<��<W��<��<��<6��<h��<1��<��<1��<��<��<��<1��<��<1��<h��<6��<��<��<W��<��<��<`   `   ���<��<��<P��<��<��<���<��<<��<��<��<��< ��<��<��<��<<��<��<���<��<��<P��<��<��<`   `   ��<��<��<��<Ѐ�<*��<)��<��<��<��<��<���<��<���<��<��<��<��<)��<*��<Ѐ�<��<��<��<`   `   ���<$��<��<ހ�<.��</��<K��<4��<��<���<��<��<��<��<��<���<��<4��<K��</��<.��<ހ�<��<$��<`   `   ��<b��<��<��<D��<��<���<6��<��<���<��<#��<��<#��<��<���<��<6��<���<��<D��<��<��<b��<`   `   ��<7��<���<��<,��<��<���<E��<!��<��<���<	��<U��<	��<���<��<!��<E��<���<��<,��<��<���<7��<`   `   ��<���<��< ��<H��<1��<.��<S��<��<��<
��<��<-��<��<
��<��<��<S��<.��<1��<H��< ��<��<���<`   `   ��<���<��<���<��<-��<��<��<��<���<���<���<���<���<���<���<��<��<��<-��<��<���<��<���<`   `   '��<
��<;��<��<���<��<���<��<"��<���<��<,��<��<,��<��<���<"��<��<���<��<���<��<;��<
��<`   `   ���<��<B��<a��<B��<(��<��<��<��<��<��<5��<7��<5��<��<��<��<��<��<(��<B��<a��<B��<��<`   `   ��<��<��<��<���<���<��<��<��<��<���<��<;��<��<���<��<��<��<��<���<���<��<��<��<`   `   +��<=��<J��<)��<	��<��< ��<��<#��<=��<��<���<��<���<��<=��<#��<��< ��<��<	��<)��<J��<=��<`   `   ���<���<(��<`��<T��<���<��<���<��<��<���<���<���<���<���<��<��<���<��<���<T��<`��<(��<���<`   `   Հ�<��<ۀ�<��<��<��<��<���<��<���<��<&��<��<&��<��<���<��<���<��<��<��<��<ۀ�<��<`   `   $��<G��<��<��<��<���<	��<��<��<"��<��<��<4��<��<��<"��<��<��<	��<���<��<��<��<G��<`   `   &��<���<��<I��<��<��<��<р�<���<��<��<��<1��<��<��<��<���<р�<��<��<��<I��<��<���<`   `   I��<��<р�<��<̀�<$��<O��<���<��<��<��<D��<;��<D��<��<��<��<���<O��<$��<̀�<��<р�<��<`   `   K��<)��<��<��<��<+��<-��<��<@��<��<)��<3��<��<3��<)��<��<@��<��<-��<+��<��<��<��<)��<`   `   ��<2��<-��< ��<��<4��<��<��<F��<݀�<��<��<���<��<��<݀�<F��<��<��<4��<��< ��<-��<2��<`   `   Ԁ�<��<)��<���<܀�<A��<��<@��<M��<���<>��<-��<,��<-��<>��<���<M��<@��<��<A��<܀�<���<)��<��<`   `   ��<��<2��<��<��</��<��<��<"��<��<
��<���<]��<���<
��<��<"��<��<��</��<��<��<2��<��<`   `   &��<���<���<!��<7��<��<̀�<��<���<��<���<ƀ�<	��<ƀ�<���<��<���<��<̀�<��<7��<!��<���<���<`   `   /��<��<���<?��<5��<���<���<��<��<��<W��<*��<��<*��<W��<��<��<��<���<���<5��<?��<���<��<`   `   ��<��<J��<%��<��<<��<5��<��<��<��<2��<'��<���<'��<2��<��<��<��<5��<<��<��<%��<J��<��<`   `   ��<��<1��<��<1��<h��<6��<��<��<W��<��<��<?��<��<��<W��<��<��<6��<h��<1��<��<1��<��<`   `    ��<��<��<��<<��<��<���<��<��<P��<��<��<���<��<��<P��<��<��<���<��<<��<��<��<��<`   `   ��<���<��<��<��<��<)��<*��<Ѐ�<��<��<��<��<��<��<��<Ѐ�<*��<)��<��<��<��<��<���<`   `   ��<��<��<���<��<4��<K��</��<.��<ހ�<��<$��<���<$��<��<ހ�<.��</��<K��<4��<��<���<��<��<`   `   ��<#��<��<���<��<6��<���<��<D��<��<��<b��<��<b��<��<��<D��<��<���<6��<��<���<��<#��<`   `   U��<	��<���<��<!��<E��<���<��<,��<��<���<7��<��<7��<���<��<,��<��<���<E��<!��<��<���<	��<`   `   -��<��<
��<��<��<S��<.��<1��<H��< ��<��<���<��<���<��< ��<H��<1��<.��<S��<��<��<
��<��<`   `   ���<���<���<���<��<��<��<-��<��<���<��<���<��<���<��<���<��<-��<��<��<��<���<���<���<`   `   ��<,��<��<���<"��<��<���<��<���<��<;��<
��<'��<
��<;��<��<���<��<���<��<"��<���<��<,��<`   `   ��<��<��<��<��<��<3��<��<��<��<��<.��<��<.��<��<��<��<��<3��<��<��<��<��<��<`   `   ��<��<1��<��<��<��<"��<��<#��<��<��<4��<��<4��<��<��<#��<��<"��<��<��<��<1��<��<`   `   ��<��<
��<��<��<��< ��<)��<*��<��<��<+��<��<+��<��<��<*��<)��< ��<��<��<��<
��<��<`   `   ��<��<��<��<)��<��<��<��<��<��<��<7��<��<7��<��<��<��<��<��<��<)��<��<��<��<`   `   ��<��<��<��<��<��<;��<��<��<��<��<��<��<��<��<��<��<��<;��<��<��<��<��<��<`   `   ��<��<��<��<��<*��<��<C��< ��<	��<��<��<��<��<��<	��< ��<C��<��<*��<��<��<��<��<`   `   ��<��<	��<��<)��<*��<��<��<��<��<��<��<��<��<��<��<��<��<��<*��<)��<��<	��<��<`   `   ��<��<��<��<��<2��<��<��<��<	��<��<��<��<��<��<	��<��<��<��<2��<��<��<��<��<`   `   $��<*��<��<��< ��<��<��<��<��<*��<��<��<��<��<��<*��<��<��<��<��< ��<��<��<*��<`   `   ��<��<��<��<!��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<!��<��<��<��<`   `   ��<��<��<��<��<��<��<*��<��<
��<��<��<��<��<��<
��<��<*��<��<��<��<��<��<��<`   `   s��<��<��<��<��<��<5��<��<��<#��<��<#��<��<#��<��<#��<��<��<5��<��<��<��<��<��<`   `   )��<��< ��<��<4��< ��<+��<��<��<-��<��<��<��<��<��<-��<��<��<+��< ��<4��<��< ��<��<`   `   ��<��<%��<��<3��<��<��<#��<��<��<��<"��<��<"��<��<��<��<#��<��<��<3��<��<%��<��<`   `   ��<��<(��<��<)��<!��<��<��<��<��<��<��<��<��<��<��<��<��<��<!��<)��<��<(��<��<`   `   ��<��<��<��<��<+��<��<��<��<��<��<��<#��<��<��<��<��<��<��<+��<��<��<��<��<`   `   1��<��<$��<)��<��<��<��<#��<��<��<��<��<G��<��<��<��<��<#��<��<��<��<)��<$��<��<`   `   ��<��<��<��<��<��<��<��<��<��<A��<
��<��<
��<A��<��<��<��<��<��<��<��<��<��<`   `   ��<��<��<0��<a��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<a��<0��<��<��<`   `   !��<-��<��<<��<9��<��<��<	��<��<��<��<��<��<��<��<��<��<	��<��<��<9��<<��<��<-��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   (��<��<��<��<��<��<��<��<��<��<	��<��<��<��<	��<��<��<��<��<��<��<��<��<��<`   `   )��<��<+��<��<��<��<��<��< ��</��<��<'��<*��<'��<��</��< ��<��<��<��<��<��<+��<��<`   `   ��<��<��<��<��<��<)��<��<��<��<��<��<��<��<��<��<��<��<)��<��<��<��<��<��<`   `   ��<.��<��<��<��<��<3��<��<��<��<��<��<��<��<��<��<��<��<3��<��<��<��<��<.��<`   `   ��<4��<��<��<#��<��<"��<��<��<��<1��<��<��<��<1��<��<��<��<"��<��<#��<��<��<4��<`   `   ��<+��<��<��<*��<)��< ��<��<��<��<
��<��<��<��<
��<��<��<��< ��<)��<*��<��<��<+��<`   `   ��<7��<��<��<��<��<��<��<)��<��<��<��<��<��<��<��<)��<��<��<��<��<��<��<7��<`   `   ��<��<��<��<��<��<;��<��<��<��<��<��<��<��<��<��<��<��<;��<��<��<��<��<��<`   `   ��<��<��<	��< ��<C��<��<*��<��<��<��<��<��<��<��<��<��<*��<��<C��< ��<	��<��<��<`   `   ��<��<��<��<��<��<��<*��<)��<��<	��<��<��<��<	��<��<)��<*��<��<��<��<��<��<��<`   `   ��<��<��<	��<��<��<��<2��<��<��<��<��<��<��<��<��<��<2��<��<��<��<	��<��<��<`   `   ��<��<��<*��<��<��<��<��< ��<��<��<*��<$��<*��<��<��< ��<��<��<��<��<*��<��<��<`   `   ��<��<��<��<��<��<��<��<!��<��<��<��<��<��<��<��<!��<��<��<��<��<��<��<��<`   `   ��<��<��<
��<��<*��<��<��<��<��<��<��<��<��<��<��<��<��<��<*��<��<
��<��<��<`   `   ��<#��<��<#��<��<��<5��<��<��<��<��<��<s��<��<��<��<��<��<5��<��<��<#��<��<#��<`   `   ��<��<��<-��<��<��<+��< ��<4��<��< ��<��<)��<��< ��<��<4��< ��<+��<��<��<-��<��<��<`   `   ��<"��<��<��<��<#��<��<��<3��<��<%��<��<��<��<%��<��<3��<��<��<#��<��<��<��<"��<`   `   ��<��<��<��<��<��<��<!��<)��<��<(��<��<��<��<(��<��<)��<!��<��<��<��<��<��<��<`   `   #��<��<��<��<��<��<��<+��<��<��<��<��<��<��<��<��<��<+��<��<��<��<��<��<��<`   `   G��<��<��<��<��<#��<��<��<��<)��<$��<��<1��<��<$��<)��<��<��<��<#��<��<��<��<��<`   `   ��<
��<A��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<A��<
��<`   `   ��<��<��<��<��<��<��<��<a��<0��<��<��<��<��<��<0��<a��<��<��<��<��<��<��<��<`   `   ��<��<��<��<��<	��<��<��<9��<<��<��<-��<!��<-��<��<<��<9��<��<��<	��<��<��<��<��<`   `   ��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<��<`   `   ��<��<	��<��<��<��<��<��<��<��<��<��<(��<��<��<��<��<��<��<��<��<��<	��<��<`   `   *��<'��<��</��< ��<��<��<��<��<��<+��<��<)��<��<+��<��<��<��<��<��< ��</��<��<'��<`   `   ��<��<��<��<��<��<)��<��<��<��<��<��<��<��<��<��<��<��<)��<��<��<��<��<��<`   `   x�<�<�~�<�~�<�<�~�<�~�<�~�<�~�<�<0�<I�<�~�<I�<0�<�<�~�<�~�<�~�<�~�<�<�~�<�~�<�<`   `   6�<�~�<�~�<�~�<;�<�~�<�~�<�~�<�~�<V�<F�<#�<�~�<#�<F�<V�<�~�<�~�<�~�<�~�<;�<�~�<�~�<�~�<`   `   	�<�~�<�~�<�~�<�<�<�<�<�~�<*�<�~�<�~�<�~�<�~�<�~�<*�<�~�<�<�<�<�<�~�<�~�<�~�<`   `   $�<�~�<�<�<�<�<�~�< �<�~�<�<�~�<�<Q�<�<�~�<�<�~�< �<�~�<�<�<�<�<�~�<`   `   �~�<�~�<�<#�<
�<�~�<�~�<�~�<�<i�< �<�~�<�<�~�< �<i�<�<�~�<�~�<�~�<
�<#�<�<�~�<`   `   *�<�<�<�~�<�~�<�<�~�<�~�<�~�<�<�~�<�~�<�~�<�~�<�~�<�<�~�<�~�<�~�<�<�~�<�~�<�<�<`   `   _�<@�<.�<�<�~�<(�<�~�<�~�<�~�<�~�<�<�<�<�<�<�~�<�~�<�~�<�~�<(�<�~�<�<.�<@�<`   `   �~�<�~�<�<.�<�~�<�~�<�~�<-�<c�<�<1�</�<�</�<1�<�<c�<-�<�~�<�~�<�~�<.�<�<�~�<`   `   �<�~�<�~�<2�<�~�<�<�<�~�<�<�~�<�~�<
�<�<
�<�~�<�~�<�<�~�<�<�<�~�<2�<�~�<�~�<`   `   m�<<�<�<4�<�~�<F�<J�<�~�<�~�<�~�<�~�<�<9�<�<�~�<�~�<�~�<�~�<J�<F�<�~�<4�<�<<�<`   `   �~�<�<�<�~�<�~�<(�<!�<�~�<=�</�<�~�<�<?�<�<�~�</�<=�<�~�<!�<(�<�~�<�~�<�<�<`   `   �~�<�~�<4�<�~�<�~�<$�<�<�~�<�<(�<�~�<�~�< �<�~�<�~�<(�<�<�~�<�<$�<�~�<�~�<4�<�~�<`   `   �~�<"�<.�<�~�<�<�~�<�<�~�<�~�<�~�< �<,�<�~�<,�< �<�~�<�~�<�~�<�<�~�<�<�~�<.�<"�<`   `   2�<�~�<�~�<�~�<"�<�~�<+�<8�<�~�<�~�<�<D�<�~�<D�<�<�~�<�~�<8�<+�<�~�<"�<�~�<�~�<�~�<`   `   L�<�~�<�~�<�<!�<�~�<�<4�<U�<1�<�~�<�<�~�<�<�~�<1�<U�<4�<�<�~�<!�<�<�~�<�~�<`   `   �<-�<%�<�~�<�~�<�~�<�~�<�~�<,�<!�<�~�<�<�~�<�<�~�<!�<,�<�~�<�~�<�~�<�~�<�~�<%�<-�<`   `   �~�<�<�<�~�<$�<%�<�<(�<�~�<�~�<�<�<�~�<�<�<�~�<�~�<(�<�<%�<$�<�~�<�<�<`   `   �~�<$�<�<�<$�<�<�<A�<�<�~�<�<�~�<�~�<�~�<�<�~�<�<A�<�<�<$�<�<�<$�<`   `   A�<�<�<�~�<�~�<�~�<�<�~�<*�<�~�<�~�<�<7�<�<�~�<�~�<*�<�~�<�<�~�<�~�<�~�<�<�<`   `   �~�<�~�<�<�~�<�~�<A�<6�<�~�<�<�<�~�<#�<�<#�<�~�<�<�<�~�<6�<A�<�~�<�~�<�<�~�<`   `   �<�~�<8�< �<�~�<R�<�<�~�<0�<�<�<&�<�~�<&�<�<�<0�<�~�<�<R�<�~�< �<8�<�~�<`   `   <�<�<�<�<�<	�<�~�<,�<<�<�~�<�~�<�<�~�<�<�~�<�~�<<�<,�<�~�<	�<�<�<�<�<`   `   
�<�<�~�<�~�<$�<�~�<�~�<:�<�<�~�<�~�<�~�<�~�<�~�<�~�<�~�<�<:�<�~�<�~�<$�<�~�<�~�<�<`   `   �~�<�<�~�<�~�<0�<!�<$�<�<�~�<�~�<�~�<�~�<%�<�~�<�~�<�~�<�~�<�<$�<!�<0�<�~�<�~�<�<`   `   �~�<I�<0�<�<�~�<�~�<�~�<�~�<�<�~�<�~�<�<x�<�<�~�<�~�<�<�~�<�~�<�~�<�~�<�<0�<I�<`   `   �~�<#�<F�<V�<�~�<�~�<�~�<�~�<;�<�~�<�~�<�~�<6�<�~�<�~�<�~�<;�<�~�<�~�<�~�<�~�<V�<F�<#�<`   `   �~�<�~�<�~�<*�<�~�<�<�<�<�<�~�<�~�<�~�<	�<�~�<�~�<�~�<�<�<�<�<�~�<*�<�~�<�~�<`   `   Q�<�<�~�<�<�~�< �<�~�<�<�<�<�<�~�<$�<�~�<�<�<�<�<�~�< �<�~�<�<�~�<�<`   `   �<�~�< �<i�<�<�~�<�~�<�~�<
�<#�<�<�~�<�~�<�~�<�<#�<
�<�~�<�~�<�~�<�<i�< �<�~�<`   `   �~�<�~�<�~�<�<�~�<�~�<�~�<�<�~�<�~�<�<�<*�<�<�<�~�<�~�<�<�~�<�~�<�~�<�<�~�<�~�<`   `   �<�<�<�~�<�~�<�~�<�~�<(�<�~�<�<.�<@�<_�<@�<.�<�<�~�<(�<�~�<�~�<�~�<�~�<�<�<`   `   �</�<1�<�<c�<-�<�~�<�~�<�~�<.�<�<�~�<�~�<�~�<�<.�<�~�<�~�<�~�<-�<c�<�<1�</�<`   `   �<
�<�~�<�~�<�<�~�<�<�<�~�<2�<�~�<�~�<�<�~�<�~�<2�<�~�<�<�<�~�<�<�~�<�~�<
�<`   `   9�<�<�~�<�~�<�~�<�~�<J�<F�<�~�<4�<�<<�<m�<<�<�<4�<�~�<F�<J�<�~�<�~�<�~�<�~�<�<`   `   ?�<�<�~�</�<=�<�~�<!�<(�<�~�<�~�<�<�<�~�<�<�<�~�<�~�<(�<!�<�~�<=�</�<�~�<�<`   `    �<�~�<�~�<(�<�<�~�<�<$�<�~�<�~�<4�<�~�<�~�<�~�<4�<�~�<�~�<$�<�<�~�<�<(�<�~�<�~�<`   `   �~�<,�< �<�~�<�~�<�~�<�<�~�<�<�~�<.�<"�<�~�<"�<.�<�~�<�<�~�<�<�~�<�~�<�~�< �<,�<`   `   �~�<D�<�<�~�<�~�<8�<+�<�~�<"�<�~�<�~�<�~�<2�<�~�<�~�<�~�<"�<�~�<+�<8�<�~�<�~�<�<D�<`   `   �~�<�<�~�<1�<U�<4�<�<�~�<!�<�<�~�<�~�<L�<�~�<�~�<�<!�<�~�<�<4�<U�<1�<�~�<�<`   `   �~�<�<�~�<!�<,�<�~�<�~�<�~�<�~�<�~�<%�<-�<�<-�<%�<�~�<�~�<�~�<�~�<�~�<,�<!�<�~�<�<`   `   �~�<�<�<�~�<�~�<(�<�<%�<$�<�~�<�<�<�~�<�<�<�~�<$�<%�<�<(�<�~�<�~�<�<�<`   `   �~�<�~�<�<�~�<�<A�<�<�<$�<�<�<$�<�~�<$�<�<�<$�<�<�<A�<�<�~�<�<�~�<`   `   7�<�<�~�<�~�<*�<�~�<�<�~�<�~�<�~�<�<�<A�<�<�<�~�<�~�<�~�<�<�~�<*�<�~�<�~�<�<`   `   �<#�<�~�<�<�<�~�<6�<A�<�~�<�~�<�<�~�<�~�<�~�<�<�~�<�~�<A�<6�<�~�<�<�<�~�<#�<`   `   �~�<&�<�<�<0�<�~�<�<R�<�~�< �<8�<�~�<�<�~�<8�< �<�~�<R�<�<�~�<0�<�<�<&�<`   `   �~�<�<�~�<�~�<<�<,�<�~�<	�<�<�<�<�<<�<�<�<�<�<	�<�~�<,�<<�<�~�<�~�<�<`   `   �~�<�~�<�~�<�~�<�<:�<�~�<�~�<$�<�~�<�~�<�<
�<�<�~�<�~�<$�<�~�<�~�<:�<�<�~�<�~�<�~�<`   `   %�<�~�<�~�<�~�<�~�<�<$�<!�<0�<�~�<�~�<�<�~�<�<�~�<�~�<0�<!�<$�<�<�~�<�~�<�~�<�~�<`   `   ,~�<�}�< ~�<~�<�}�<~�<~�<c~�<�}�<�}�<�}�<�}�<	~�<�}�<�}�<�}�<�}�<c~�<~�<~�<�}�<~�< ~�<�}�<`   `   ~�<�}�<5~�<'~�<~�<~�<~�<J~�<�}�<	~�<�}�<�}�<V~�<�}�<�}�<	~�<�}�<J~�<~�<~�<~�<'~�<5~�<�}�<`   `   ~�< ~�<F~�<#~�<�}�<#~�<�}�<
~�<�}�<~�<~�<~�<s~�<~�<~�<~�<�}�<
~�<�}�<#~�<�}�<#~�<F~�< ~�<`   `   G~�<~�<~�< ~�<�}�<5~�<~�<0~�<7~�<�}�<.~�<~�<�}�<~�<.~�<�}�<7~�<0~�<~�<5~�<�}�< ~�<~�<~�<`   `   3~�<~�<�}�<*~�<+~�<-~�<~�<7~�<$~�<�}�<~�<	~�<�}�<	~�<~�<�}�<$~�<7~�<~�<-~�<+~�<*~�<�}�<~�<`   `   �}�<~�<�}�<"~�<&~�<�}�<6~�<~�<~�<~�<~�<=~�<n~�<=~�<~�<~�<~�<~�<6~�<�}�<&~�<"~�<�}�<~�<`   `   �}�<~�<�}�<~�<&~�<~�<l~�<~�<~�<@~�<
~�<~�<)~�<~�<
~�<@~�<~�<~�<l~�<~�<&~�<~�<�}�<~�<`   `   -~�<L~�<~�<&~�<H~�<�}�<~�<�}�<�}�<~�<�}�<�}�<�}�<�}�<�}�<~�<�}�<�}�<~�<�}�<H~�<&~�<~�<L~�<`   `   �}�<+~�<~�<~�<~�<�}�<�}�<~�<	~�<~�<~�< ~�<~�< ~�<~�<~�<	~�<~�<�}�<�}�<~�<~�<~�<+~�<`   `   �}�<~�<~�<�}�<	~�<~�<~�<=~�<%~�<7~�<p~�<�}�<�}�<�}�<p~�<7~�<%~�<=~�<~�<~�<	~�<�}�<~�<~�<`   `   3~�<;~�<�}�<)~�<6~�<�}�<�}�<%~�<�}�<�}�<j~�<�}�<�}�<�}�<j~�<�}�<�}�<%~�<�}�<�}�<6~�<)~�<�}�<;~�<`   `   ;~�<)~�<�}�<~�<E~�<~�<�}�<q~�<*~�<�}�<'~�<~�<~�<~�<'~�<�}�<*~�<q~�<�}�<~�<E~�<~�<�}�<)~�<`   `   7~�<0~�<#~�<	~�<~�<!~�<�}�<6~�<:~�<+~�<%~�<~�<.~�<~�<%~�<+~�<:~�<6~�<�}�<!~�<~�<	~�<#~�<0~�<`   `   ~�<�}�<>~�<+~�<�}�<~�<�}�<�}�<�}�</~�<�}�<�}�<~�<�}�<�}�</~�<�}�<�}�<�}�<~�<�}�<+~�<>~�<�}�<`   `   �}�<�}�<=~�<V~�<~�<)~�<J~�<�}�<�}�<~�<�}�<~�<&~�<~�<�}�<~�<�}�<�}�<J~�<)~�<~�<V~�<=~�<�}�<`   `   &~�<!~�<6~�<O~�< ~�<~�<B~�<~�<�}�<	~�<~�<E~�<,~�<E~�<~�<	~�<�}�<~�<B~�<~�< ~�<O~�<6~�<!~�<`   `   ~�<~�<�}�<~�<.~�<�}�< ~�<�}�<~�<~�<~�<~�<�}�<~�<~�<~�<~�<�}�< ~�<�}�<.~�<~�<�}�<~�<`   `   ~�<~�<~�<,~�<~�<~�<�}�<�}�<;~�<6~�<~�<~�<~�<~�<~�<6~�<;~�<�}�<�}�<~�<~�<,~�<~�<~�<`   `   ~�<�}�<'~�<L~�<3~�<>~�<~�<�}�<�}�<~�<9~�<~�<~�<~�<9~�<~�<�}�<�}�<~�<>~�<3~�<L~�<'~�<�}�<`   `   B~�<!~�<~�<-~�<[~�<~�<�}�<9~�<�}�<�}�<~�<�}�<�}�<�}�<~�<�}�<�}�<9~�<�}�<~�<[~�<-~�<~�<!~�<`   `   U~�<M~�<~�<~�<G~�<�}�<�}�<;~�<~�<~�<�}�<~�<~�<~�<�}�<~�<~�<;~�<�}�<�}�<G~�<~�<~�<M~�<`   `   �}�<�}�< ~�<�}�<~�<~�</~�<~�<�}�<~�<~�<3~�<0~�<3~�<~�<~�<�}�<~�</~�<~�<~�<�}�< ~�<�}�<`   `   ~�<~�<)~�<~�<�}�<~�<#~�<�}�<�}�<A~�<G~�<~�<�}�<~�<G~�<A~�<�}�<�}�<#~�<~�<�}�<~�<)~�<~�<`   `   <~�<4~�<5~�<'~�<~�<	~�<�}�<~�<~�<3~�<L~�<�}�<�}�<�}�<L~�<3~�<~�<~�<�}�<	~�<~�<'~�<5~�<4~�<`   `   	~�<�}�<�}�<�}�<�}�<c~�<~�<~�<�}�<~�< ~�<�}�<,~�<�}�< ~�<~�<�}�<~�<~�<c~�<�}�<�}�<�}�<�}�<`   `   V~�<�}�<�}�<	~�<�}�<J~�<~�<~�<~�<'~�<5~�<�}�<~�<�}�<5~�<'~�<~�<~�<~�<J~�<�}�<	~�<�}�<�}�<`   `   s~�<~�<~�<~�<�}�<
~�<�}�<#~�<�}�<#~�<F~�< ~�<~�< ~�<F~�<#~�<�}�<#~�<�}�<
~�<�}�<~�<~�<~�<`   `   �}�<~�<.~�<�}�<7~�<0~�<~�<5~�<�}�< ~�<~�<~�<G~�<~�<~�< ~�<�}�<5~�<~�<0~�<7~�<�}�<.~�<~�<`   `   �}�<	~�<~�<�}�<$~�<7~�<~�<-~�<+~�<*~�<�}�<~�<3~�<~�<�}�<*~�<+~�<-~�<~�<7~�<$~�<�}�<~�<	~�<`   `   n~�<=~�<~�<~�<~�<~�<6~�<�}�<&~�<"~�<�}�<~�<�}�<~�<�}�<"~�<&~�<�}�<6~�<~�<~�<~�<~�<=~�<`   `   )~�<~�<
~�<@~�<~�<~�<l~�<~�<&~�<~�<�}�<~�<�}�<~�<�}�<~�<&~�<~�<l~�<~�<~�<@~�<
~�<~�<`   `   �}�<�}�<�}�<~�<�}�<�}�<~�<�}�<H~�<&~�<~�<L~�<-~�<L~�<~�<&~�<H~�<�}�<~�<�}�<�}�<~�<�}�<�}�<`   `   ~�< ~�<~�<~�<	~�<~�<�}�<�}�<~�<~�<~�<+~�<�}�<+~�<~�<~�<~�<�}�<�}�<~�<	~�<~�<~�< ~�<`   `   �}�<�}�<p~�<7~�<%~�<=~�<~�<~�<	~�<�}�<~�<~�<�}�<~�<~�<�}�<	~�<~�<~�<=~�<%~�<7~�<p~�<�}�<`   `   �}�<�}�<j~�<�}�<�}�<%~�<�}�<�}�<6~�<)~�<�}�<;~�<3~�<;~�<�}�<)~�<6~�<�}�<�}�<%~�<�}�<�}�<j~�<�}�<`   `   ~�<~�<'~�<�}�<*~�<q~�<�}�<~�<E~�<~�<�}�<)~�<;~�<)~�<�}�<~�<E~�<~�<�}�<q~�<*~�<�}�<'~�<~�<`   `   .~�<~�<%~�<+~�<:~�<6~�<�}�<!~�<~�<	~�<#~�<0~�<7~�<0~�<#~�<	~�<~�<!~�<�}�<6~�<:~�<+~�<%~�<~�<`   `   ~�<�}�<�}�</~�<�}�<�}�<�}�<~�<�}�<+~�<>~�<�}�<~�<�}�<>~�<+~�<�}�<~�<�}�<�}�<�}�</~�<�}�<�}�<`   `   &~�<~�<�}�<~�<�}�<�}�<J~�<)~�<~�<V~�<=~�<�}�<�}�<�}�<=~�<V~�<~�<)~�<J~�<�}�<�}�<~�<�}�<~�<`   `   ,~�<E~�<~�<	~�<�}�<~�<B~�<~�< ~�<O~�<6~�<!~�<&~�<!~�<6~�<O~�< ~�<~�<B~�<~�<�}�<	~�<~�<E~�<`   `   �}�<~�<~�<~�<~�<�}�< ~�<�}�<.~�<~�<�}�<~�<~�<~�<�}�<~�<.~�<�}�< ~�<�}�<~�<~�<~�<~�<`   `   ~�<~�<~�<6~�<;~�<�}�<�}�<~�<~�<,~�<~�<~�<~�<~�<~�<,~�<~�<~�<�}�<�}�<;~�<6~�<~�<~�<`   `   ~�<~�<9~�<~�<�}�<�}�<~�<>~�<3~�<L~�<'~�<�}�<~�<�}�<'~�<L~�<3~�<>~�<~�<�}�<�}�<~�<9~�<~�<`   `   �}�<�}�<~�<�}�<�}�<9~�<�}�<~�<[~�<-~�<~�<!~�<B~�<!~�<~�<-~�<[~�<~�<�}�<9~�<�}�<�}�<~�<�}�<`   `   ~�<~�<�}�<~�<~�<;~�<�}�<�}�<G~�<~�<~�<M~�<U~�<M~�<~�<~�<G~�<�}�<�}�<;~�<~�<~�<�}�<~�<`   `   0~�<3~�<~�<~�<�}�<~�</~�<~�<~�<�}�< ~�<�}�<�}�<�}�< ~�<�}�<~�<~�</~�<~�<�}�<~�<~�<3~�<`   `   �}�<~�<G~�<A~�<�}�<�}�<#~�<~�<�}�<~�<)~�<~�<~�<~�<)~�<~�<�}�<~�<#~�<�}�<�}�<A~�<G~�<~�<`   `   �}�<�}�<L~�<3~�<~�<~�<�}�<	~�<~�<'~�<5~�<4~�<<~�<4~�<5~�<'~�<~�<	~�<�}�<~�<~�<3~�<L~�<�}�<`   `   }�<0}�<?}�<}�<&}�<T}�<$}�<}�<@}�<F}�<C}�</}�<6}�</}�<C}�<F}�<@}�<}�<$}�<T}�<&}�<}�<?}�<0}�<`   `   (}�<U}�<}�<}�< }�<'}�<2}�<$}�<>}�<8}�<H}�<<}�<L}�<<}�<H}�<8}�<>}�<$}�<2}�<'}�< }�<}�<}�<U}�<`   `   &}�<T}�<}�<T}�<V}�<,}�<$}�<}�<O}�<%}�<>}�<'}�<(}�<'}�<>}�<%}�<O}�<}�<$}�<,}�<V}�<T}�<}�<T}�<`   `   �|�<#}�<}�<8}�<}�<5}�<*}�<}�<S}�<}�<`}�</}�<}�</}�<`}�<}�<S}�<}�<*}�<5}�<}�<8}�<}�<#}�<`   `   !}�<[}�<$}�<}�<}�<F}�<2}�<}�<,}�<�|�<F}�<<}�<#}�<<}�<F}�<�|�<,}�<}�<2}�<F}�<}�<}�<$}�<[}�<`   `   <}�<u}�<_}�<M}�<?}�<}�<
}�<}�<J}�<:}�<*}�<,}�<}�<,}�<*}�<:}�<J}�<}�<
}�<}�<?}�<M}�<_}�<u}�<`   `   �|�<}�<7}�<(}�<%}�<�|�<%}�<#}�<T}�<e}�</}�<#}�<�|�<#}�</}�<e}�<T}�<#}�<%}�<�|�<%}�<(}�<7}�<}�<`   `   =}�<B}�<0}�<}�<<}�<3}�<A}�<}�<}�<)}�<0}�<]}�<4}�<]}�<0}�<)}�<}�<}�<A}�<3}�<<}�<}�<0}�<B}�<`   `   C}�<U}�<L}�<}�<J}�<@}�</}�<L}�<1}�<9}�<}�<Q}�<�}�<Q}�<}�<9}�<1}�<L}�</}�<@}�<J}�<}�<L}�<U}�<`   `   �|�<}�<A}�<"}�<*}�<C}�<2}�<O}�<K}�<:}�<�|�<�|�<^}�<�|�<�|�<:}�<K}�<O}�<2}�<C}�<*}�<"}�<A}�<}�<`   `   ?}�<D}�<A}�<V}�<}�<=}�<9}�<}�<}�<}�<}�<}�<s}�<}�<}�<}�<}�<}�<9}�<=}�<}�<V}�<A}�<D}�<`   `   2}�<}�<}�<O}�<�|�<&}�<N}�<%}�<}�<0}�<T}�<*}�<s}�<*}�<T}�<0}�<}�<%}�<N}�<&}�<�|�<O}�<}�<}�<`   `   }�<
}�<}�<?}�<}�<S}�<F}�<7}�<$}�<8}�<8}�<�|�<Z}�<�|�<8}�<8}�<$}�<7}�<F}�<S}�<}�<?}�<}�<
}�<`   `   V}�<S}�<E}�<}�<4}�<t}�<}�<H}�<<}�<-}�<9}�<}�<l}�<}�<9}�<-}�<<}�<H}�<}�<t}�<4}�<}�<E}�<S}�<`   `   V}�<A}�<}�<�|�<}�<3}�<�|�<P}�<9}�<"}�<R}�<"}�<'}�<"}�<R}�<"}�<9}�<P}�<�|�<3}�<}�<�|�<}�<A}�<`   `   ,}�</}�<}�<}�<;}�<'}�<+}�<9}�<*}�<9}�<I}�<}�<�|�<}�<I}�<9}�<*}�<9}�<+}�<'}�<;}�<}�<}�</}�<`   `   8}�<E}�<,}�<@}�<5}�<>}�<j}�<:}�<J}�<A}�<}�<$}�<G}�<$}�<}�<A}�<J}�<:}�<j}�<>}�<5}�<@}�<,}�<E}�<`   `   C}�<D}�<=}�<}�<�|�<1}�<P}�<%}�<+}�<}�<}�<8}�<_}�<8}�<}�<}�<+}�<%}�<P}�<1}�<�|�<}�<=}�<D}�<`   `   }�<*}�<:}�<}�<!}�<>}�<:}�<K}�<}�<'}�<J}�<&}�<*}�<&}�<J}�<'}�<}�<K}�<:}�<>}�<!}�<}�<:}�<*}�<`   `   �|�<0}�<}�<�|�<G}�<
}�<0}�<u}�<"}�<I}�<9}�<}�<V}�<}�<9}�<I}�<"}�<u}�<0}�<
}�<G}�<�|�<}�<0}�<`   `   �|�<@}�<%}�<	}�<-}�<�|�<R}�<5}�<}�<^}�<%}�<)}�<Y}�<)}�<%}�<^}�<}�<5}�<R}�<�|�<-}�<	}�<%}�<@}�<`   `   }�<,}�<B}�<O}�<2}�<S}�<�}�<�|�< }�<]}�<}�<}�<}�<}�<}�<]}�< }�<�|�<�}�<S}�<2}�<O}�<B}�<,}�<`   `   O}�<-}�<-}�<M}�<%}�<G}�<I}�<}�<L}�<}�<�|�<5}�<I}�<5}�<�|�<}�<L}�<}�<I}�<G}�<%}�<M}�<-}�<-}�<`   `   P}�<'}�<}�<5}�<*}�<}�<}�<i}�<e}�<}�<}�<?}�<b}�<?}�<}�<}�<e}�<i}�<}�<}�<*}�<5}�<}�<'}�<`   `   6}�</}�<C}�<F}�<@}�<}�<$}�<T}�<&}�<}�<?}�<0}�<}�<0}�<?}�<}�<&}�<T}�<$}�<}�<@}�<F}�<C}�</}�<`   `   L}�<<}�<H}�<8}�<>}�<$}�<2}�<'}�< }�<}�<}�<U}�<(}�<U}�<}�<}�< }�<'}�<2}�<$}�<>}�<8}�<H}�<<}�<`   `   (}�<'}�<>}�<%}�<O}�<}�<$}�<,}�<V}�<T}�<}�<T}�<&}�<T}�<}�<T}�<V}�<,}�<$}�<}�<O}�<%}�<>}�<'}�<`   `   }�</}�<`}�<}�<S}�<}�<*}�<5}�<}�<8}�<}�<#}�<�|�<#}�<}�<8}�<}�<5}�<*}�<}�<S}�<}�<`}�</}�<`   `   #}�<<}�<F}�<�|�<,}�<}�<2}�<F}�<}�<}�<$}�<[}�<!}�<[}�<$}�<}�<}�<F}�<2}�<}�<,}�<�|�<F}�<<}�<`   `   }�<,}�<*}�<:}�<J}�<}�<
}�<}�<?}�<M}�<_}�<u}�<<}�<u}�<_}�<M}�<?}�<}�<
}�<}�<J}�<:}�<*}�<,}�<`   `   �|�<#}�</}�<e}�<T}�<#}�<%}�<�|�<%}�<(}�<7}�<}�<�|�<}�<7}�<(}�<%}�<�|�<%}�<#}�<T}�<e}�</}�<#}�<`   `   4}�<]}�<0}�<)}�<}�<}�<A}�<3}�<<}�<}�<0}�<B}�<=}�<B}�<0}�<}�<<}�<3}�<A}�<}�<}�<)}�<0}�<]}�<`   `   �}�<Q}�<}�<9}�<1}�<L}�</}�<@}�<J}�<}�<L}�<U}�<C}�<U}�<L}�<}�<J}�<@}�</}�<L}�<1}�<9}�<}�<Q}�<`   `   ^}�<�|�<�|�<:}�<K}�<O}�<2}�<C}�<*}�<"}�<A}�<}�<�|�<}�<A}�<"}�<*}�<C}�<2}�<O}�<K}�<:}�<�|�<�|�<`   `   s}�<}�<}�<}�<}�<}�<9}�<=}�<}�<V}�<A}�<D}�<?}�<D}�<A}�<V}�<}�<=}�<9}�<}�<}�<}�<}�<}�<`   `   s}�<*}�<T}�<0}�<}�<%}�<N}�<&}�<�|�<O}�<}�<}�<2}�<}�<}�<O}�<�|�<&}�<N}�<%}�<}�<0}�<T}�<*}�<`   `   Z}�<�|�<8}�<8}�<$}�<7}�<F}�<S}�<}�<?}�<}�<
}�<}�<
}�<}�<?}�<}�<S}�<F}�<7}�<$}�<8}�<8}�<�|�<`   `   l}�<}�<9}�<-}�<<}�<H}�<}�<t}�<4}�<}�<E}�<S}�<V}�<S}�<E}�<}�<4}�<t}�<}�<H}�<<}�<-}�<9}�<}�<`   `   '}�<"}�<R}�<"}�<9}�<P}�<�|�<3}�<}�<�|�<}�<A}�<V}�<A}�<}�<�|�<}�<3}�<�|�<P}�<9}�<"}�<R}�<"}�<`   `   �|�<}�<I}�<9}�<*}�<9}�<+}�<'}�<;}�<}�<}�</}�<,}�</}�<}�<}�<;}�<'}�<+}�<9}�<*}�<9}�<I}�<}�<`   `   G}�<$}�<}�<A}�<J}�<:}�<j}�<>}�<5}�<@}�<,}�<E}�<8}�<E}�<,}�<@}�<5}�<>}�<j}�<:}�<J}�<A}�<}�<$}�<`   `   _}�<8}�<}�<}�<+}�<%}�<P}�<1}�<�|�<}�<=}�<D}�<C}�<D}�<=}�<}�<�|�<1}�<P}�<%}�<+}�<}�<}�<8}�<`   `   *}�<&}�<J}�<'}�<}�<K}�<:}�<>}�<!}�<}�<:}�<*}�<}�<*}�<:}�<}�<!}�<>}�<:}�<K}�<}�<'}�<J}�<&}�<`   `   V}�<}�<9}�<I}�<"}�<u}�<0}�<
}�<G}�<�|�<}�<0}�<�|�<0}�<}�<�|�<G}�<
}�<0}�<u}�<"}�<I}�<9}�<}�<`   `   Y}�<)}�<%}�<^}�<}�<5}�<R}�<�|�<-}�<	}�<%}�<@}�<�|�<@}�<%}�<	}�<-}�<�|�<R}�<5}�<}�<^}�<%}�<)}�<`   `   }�<}�<}�<]}�< }�<�|�<�}�<S}�<2}�<O}�<B}�<,}�<}�<,}�<B}�<O}�<2}�<S}�<�}�<�|�< }�<]}�<}�<}�<`   `   I}�<5}�<�|�<}�<L}�<}�<I}�<G}�<%}�<M}�<-}�<-}�<O}�<-}�<-}�<M}�<%}�<G}�<I}�<}�<L}�<}�<�|�<5}�<`   `   b}�<?}�<}�<}�<e}�<i}�<}�<}�<*}�<5}�<}�<'}�<P}�<'}�<}�<5}�<*}�<}�<}�<i}�<e}�<}�<}�<?}�<`   `   0|�<Z|�<||�<�|�<G|�<0|�<b|�</|�<_|�<M|�<y|�<�|�<8|�<�|�<y|�<M|�<_|�</|�<b|�<0|�<G|�<�|�<||�<Z|�<`   `   0|�<{|�<"|�<U|�<_|�<7|�<l|�<2|�<i|�<@|�<l|�<m|�<|�<m|�<l|�<@|�<i|�<2|�<l|�<7|�<_|�<U|�<"|�<{|�<`   `   A|�<�|�<|�<[|�<s|�<@|�<�|�<e|�<d|�<,|�<8|�<<|�<+|�<<|�<8|�<,|�<d|�<e|�<�|�<@|�<s|�<[|�<|�<�|�<`   `   7|�<�|�<x|�<�|�<U|�<&|�<o|�<E|�<Q|�<k|�<@|�<K|�<�|�<K|�<@|�<k|�<Q|�<E|�<o|�<&|�<U|�<�|�<x|�<�|�<`   `   "|�<2|�<=|�<R|�<;|�<S|�<t|�<d|�<\|�<�|�<T|�<2|�<�|�<2|�<T|�<�|�<\|�<d|�<t|�<S|�<;|�<R|�<=|�<2|�<`   `   �|�<4|�<*|�<6|�<a|�<�|�<c|�<o|�<E|�<R|�<V|�<@|�<W|�<@|�<V|�<R|�<E|�<o|�<c|�<�|�<a|�<6|�<*|�<4|�<`   `   �|�<J|�<v|�<V|�<R|�<�|�<G|�<b|�<A|�<|�<<|�<�|�<i|�<�|�<<|�<|�<A|�<b|�<G|�<�|�<R|�<V|�<v|�<J|�<`   `   a|�<�{�<r|�<c|�<7|�<m|�<[|�<�|�<u|�<E|�<I|�<s|�<+|�<s|�<I|�<E|�<u|�<�|�<[|�<m|�<7|�<c|�<r|�<�{�<`   `   �|�<|�<]|�<�|�<P|�<>|�<:|�<\|�<I|�<n|�<v|�<K|�<�{�<K|�<v|�<n|�<I|�<\|�<:|�<>|�<P|�<�|�<]|�<|�<`   `   �|�<J|�<E|�<b|�<V|�<W|�<K|�<)|�<&|�<E|�<Z|�<s|�<<|�<s|�<Z|�<E|�<&|�<)|�<K|�<W|�<V|�<b|�<E|�<J|�<`   `   L|�<T|�<P|�<D|�<L|�<�|�<�|�<B|�<�|�<�|�<L|�<||�<c|�<||�<L|�<�|�<�|�<B|�<�|�<�|�<L|�<D|�<P|�<T|�<`   `   2|�<�|�<r|�<b|�<M|�<T|�<V|�<|�<�|�<�|�<P|�<F|�<|�<F|�<P|�<�|�<�|�<|�<V|�<T|�<M|�<b|�<r|�<�|�<`   `   C|�<y|�<P|�<o|�<U|�<|�<>|�<%|�<-|�<%|�<Q|�<J|�<.|�<J|�<Q|�<%|�<-|�<%|�<>|�<|�<U|�<o|�<P|�<y|�<`   `   =|�<W|�<J|�<�|�<o|�<8|�<]|�<�|�<a|�<9|�<~|�<i|�<_|�<i|�<~|�<9|�<a|�<�|�<]|�<8|�<o|�<�|�<J|�<W|�<`   `   <|�<`|�<t|�<�|�<�|�<S|�<;|�<{|�<k|�<D|�<l|�<U|�<Z|�<U|�<l|�<D|�<k|�<{|�<;|�<S|�<�|�<�|�<t|�<`|�<`   `   .|�<k|�<�|�<m|�<i|�<V|�<2|�<B|�<M|�<I|�<L|�<P|�<p|�<P|�<L|�<I|�<M|�<B|�<2|�<V|�<i|�<m|�<�|�<k|�<`   `    |�<R|�<p|�<c|�<a|�<Z|�<M|�<K|�<U|�<d|�<m|�<h|�<j|�<h|�<m|�<d|�<U|�<K|�<M|�<Z|�<a|�<c|�<p|�<R|�<`   `   M|�<<|�<G|�<m|�<w|�<b|�<>|�<S|�<P|�<<|�<p|�<[|�<%|�<[|�<p|�<<|�<P|�<S|�<>|�<b|�<w|�<m|�<G|�<<|�<`   `   �|�<g|�<\|�<i|�<[|�<^|�<-|�<P|�<�|�<Y|�<S|�<D|�<(|�<D|�<S|�<Y|�<�|�<P|�<-|�<^|�<[|�<i|�<\|�<g|�<`   `   u|�<h|�<z|�<l|�<G|�<�|�<S|�<|�<c|�<`|�<2|�<\|�<�|�<\|�<2|�<`|�<c|�<|�<S|�<�|�<G|�<l|�<z|�<h|�<`   `   ]|�<O|�<a|�<|�<[|�<�|�<o|�<(|�<T|�<4|�<D|�<m|�<\|�<m|�<D|�<4|�<T|�<(|�<o|�<�|�<[|�<|�<a|�<O|�<`   `   �|�<p|�<P|�<p|�<H|�<'|�<|�<t|�<�|�<@|�<�|�<r|�<�{�<r|�<�|�<@|�<�|�<t|�<|�<'|�<H|�<p|�<P|�<p|�<`   `   `|�<W|�<=|�<?|�<W|�<M|�<|�<W|�<m|�<&|�<e|�<s|�<D|�<s|�<e|�<&|�<m|�<W|�<|�<M|�<W|�<?|�<=|�<W|�<`   `   |�<A|�<A|�<0|�<s|�<�|�<~|�<:|�<#|�<^|�<Y|�<O|�<c|�<O|�<Y|�<^|�<#|�<:|�<~|�<�|�<s|�<0|�<A|�<A|�<`   `   8|�<�|�<y|�<M|�<_|�</|�<b|�<0|�<G|�<�|�<||�<Z|�<0|�<Z|�<||�<�|�<G|�<0|�<b|�</|�<_|�<M|�<y|�<�|�<`   `   |�<m|�<l|�<@|�<i|�<2|�<l|�<7|�<_|�<U|�<"|�<{|�<0|�<{|�<"|�<U|�<_|�<7|�<l|�<2|�<i|�<@|�<l|�<m|�<`   `   +|�<<|�<8|�<,|�<d|�<e|�<�|�<@|�<s|�<[|�<|�<�|�<A|�<�|�<|�<[|�<s|�<@|�<�|�<e|�<d|�<,|�<8|�<<|�<`   `   �|�<K|�<@|�<k|�<Q|�<E|�<o|�<&|�<U|�<�|�<x|�<�|�<7|�<�|�<x|�<�|�<U|�<&|�<o|�<E|�<Q|�<k|�<@|�<K|�<`   `   �|�<2|�<T|�<�|�<\|�<d|�<t|�<S|�<;|�<R|�<=|�<2|�<"|�<2|�<=|�<R|�<;|�<S|�<t|�<d|�<\|�<�|�<T|�<2|�<`   `   W|�<@|�<V|�<R|�<E|�<o|�<c|�<�|�<a|�<6|�<*|�<4|�<�|�<4|�<*|�<6|�<a|�<�|�<c|�<o|�<E|�<R|�<V|�<@|�<`   `   i|�<�|�<<|�<|�<A|�<b|�<G|�<�|�<R|�<V|�<v|�<J|�<�|�<J|�<v|�<V|�<R|�<�|�<G|�<b|�<A|�<|�<<|�<�|�<`   `   +|�<s|�<I|�<E|�<u|�<�|�<[|�<m|�<7|�<c|�<r|�<�{�<a|�<�{�<r|�<c|�<7|�<m|�<[|�<�|�<u|�<E|�<I|�<s|�<`   `   �{�<K|�<v|�<n|�<I|�<\|�<:|�<>|�<P|�<�|�<]|�<|�<�|�<|�<]|�<�|�<P|�<>|�<:|�<\|�<I|�<n|�<v|�<K|�<`   `   <|�<s|�<Z|�<E|�<&|�<)|�<K|�<W|�<V|�<b|�<E|�<J|�<�|�<J|�<E|�<b|�<V|�<W|�<K|�<)|�<&|�<E|�<Z|�<s|�<`   `   c|�<||�<L|�<�|�<�|�<B|�<�|�<�|�<L|�<D|�<P|�<T|�<L|�<T|�<P|�<D|�<L|�<�|�<�|�<B|�<�|�<�|�<L|�<||�<`   `   |�<F|�<P|�<�|�<�|�<|�<V|�<T|�<M|�<b|�<r|�<�|�<2|�<�|�<r|�<b|�<M|�<T|�<V|�<|�<�|�<�|�<P|�<F|�<`   `   .|�<J|�<Q|�<%|�<-|�<%|�<>|�<|�<U|�<o|�<P|�<y|�<C|�<y|�<P|�<o|�<U|�<|�<>|�<%|�<-|�<%|�<Q|�<J|�<`   `   _|�<i|�<~|�<9|�<a|�<�|�<]|�<8|�<o|�<�|�<J|�<W|�<=|�<W|�<J|�<�|�<o|�<8|�<]|�<�|�<a|�<9|�<~|�<i|�<`   `   Z|�<U|�<l|�<D|�<k|�<{|�<;|�<S|�<�|�<�|�<t|�<`|�<<|�<`|�<t|�<�|�<�|�<S|�<;|�<{|�<k|�<D|�<l|�<U|�<`   `   p|�<P|�<L|�<I|�<M|�<B|�<2|�<V|�<i|�<m|�<�|�<k|�<.|�<k|�<�|�<m|�<i|�<V|�<2|�<B|�<M|�<I|�<L|�<P|�<`   `   j|�<h|�<m|�<d|�<U|�<K|�<M|�<Z|�<a|�<c|�<p|�<R|�< |�<R|�<p|�<c|�<a|�<Z|�<M|�<K|�<U|�<d|�<m|�<h|�<`   `   %|�<[|�<p|�<<|�<P|�<S|�<>|�<b|�<w|�<m|�<G|�<<|�<M|�<<|�<G|�<m|�<w|�<b|�<>|�<S|�<P|�<<|�<p|�<[|�<`   `   (|�<D|�<S|�<Y|�<�|�<P|�<-|�<^|�<[|�<i|�<\|�<g|�<�|�<g|�<\|�<i|�<[|�<^|�<-|�<P|�<�|�<Y|�<S|�<D|�<`   `   �|�<\|�<2|�<`|�<c|�<|�<S|�<�|�<G|�<l|�<z|�<h|�<u|�<h|�<z|�<l|�<G|�<�|�<S|�<|�<c|�<`|�<2|�<\|�<`   `   \|�<m|�<D|�<4|�<T|�<(|�<o|�<�|�<[|�<|�<a|�<O|�<]|�<O|�<a|�<|�<[|�<�|�<o|�<(|�<T|�<4|�<D|�<m|�<`   `   �{�<r|�<�|�<@|�<�|�<t|�<|�<'|�<H|�<p|�<P|�<p|�<�|�<p|�<P|�<p|�<H|�<'|�<|�<t|�<�|�<@|�<�|�<r|�<`   `   D|�<s|�<e|�<&|�<m|�<W|�<|�<M|�<W|�<?|�<=|�<W|�<`|�<W|�<=|�<?|�<W|�<M|�<|�<W|�<m|�<&|�<e|�<s|�<`   `   c|�<O|�<Y|�<^|�<#|�<:|�<~|�<�|�<s|�<0|�<A|�<A|�<|�<A|�<A|�<0|�<s|�<�|�<~|�<:|�<#|�<^|�<Y|�<O|�<`   `   �{�<�{�<Z{�<�{�<�{�<�{�<�{�<u{�<�{�<�{�<M{�<y{�<�{�<y{�<M{�<�{�<�{�<u{�<�{�<�{�<�{�<�{�<Z{�<�{�<`   `   y{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<b{�<�{�<�{�<�{�<b{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<`   `   H{�<e{�<�{�<f{�<f{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<f{�<f{�<�{�<e{�<`   `   �{�<�{�<�{�<j{�<�{�<�{�<k{�<�{�<n{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<n{�<�{�<k{�<�{�<�{�<j{�<�{�<�{�<`   `   �{�<�{�<�{�<�{�<�{�<�{�<i{�<�{�<w{�<~{�<�{�<g{�<w{�<g{�<�{�<~{�<w{�<�{�<i{�<�{�<�{�<�{�<�{�<�{�<`   `   k{�<Z{�<�{�<�{�<�{�<p{�<v{�<�{�<v{�<�{�<�{�<�{�<{{�<�{�<�{�<�{�<v{�<�{�<v{�<p{�<�{�<�{�<�{�<Z{�<`   `   �{�<�{�<�{�<�{�<�{�<�{�<k{�<}{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<}{�<k{�<�{�<�{�<�{�<�{�<�{�<`   `   �{�<�{�<�{�<r{�<�{�<�{�<z{�<n{�<�{�<�{�<^{�<p{�<�{�<p{�<^{�<�{�<�{�<n{�<z{�<�{�<�{�<r{�<�{�<�{�<`   `   �{�<�{�<�{�<t{�<�{�<�{�<�{�<�{�<�{�<�{�<|{�<�{�<�{�<�{�<|{�<�{�<�{�<�{�<�{�<�{�<�{�<t{�<�{�<�{�<`   `   �{�<�{�<�{�<�{�<�{�<h{�<�{�<�{�<x{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<x{�<�{�<�{�<h{�<�{�<�{�<�{�<�{�<`   `   R{�<q{�<�{�<x{�<�{�<K{�<q{�<�{�<|{�<R{�<z{�<�{�<9{�<�{�<z{�<R{�<|{�<�{�<q{�<K{�<�{�<x{�<�{�<q{�<`   `   �{�<�{�<�{�<z{�<�{�<�{�<�{�<�{�<�{�<N{�<x{�<�{�<s{�<�{�<x{�<N{�<�{�<�{�<�{�<�{�<�{�<z{�<�{�<�{�<`   `   �{�<�{�<k{�<g{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<g{�<k{�<�{�<`   `   �{�<�{�<n{�<q{�<Z{�<�{�<�{�<S{�<�{�<�{�<{{�<v{�<l{�<v{�<{{�<�{�<�{�<S{�<�{�<�{�<Z{�<q{�<n{�<�{�<`   `   �{�<{{�<�{�<�{�<d{�<�{�<�{�<7{�<k{�<�{�<m{�<{{�<�{�<{{�<m{�<�{�<k{�<7{�<�{�<�{�<d{�<�{�<�{�<{{�<`   `   �{�<�{�<h{�<q{�<e{�<�{�<�{�<�{�<�{�<�{�<r{�<�{�<�{�<�{�<r{�<�{�<�{�<�{�<�{�<�{�<e{�<q{�<h{�<�{�<`   `   �{�<�{�<~{�<a{�<j{�<p{�<�{�<�{�<�{�<�{�<�{�<u{�<n{�<u{�<�{�<�{�<�{�<�{�<�{�<p{�<j{�<a{�<~{�<�{�<`   `   �{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<w{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<w{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<`   `   �{�<s{�<x{�<�{�<�{�<�{�<�{�<�{�<�{�<~{�<�{�<�{�<�{�<�{�<�{�<~{�<�{�<�{�<�{�<�{�<�{�<�{�<x{�<s{�<`   `   �{�<w{�<�{�<�{�<^{�<w{�<�{�<�{�<�{�<�{�<�{�<�{�<^{�<�{�<�{�<�{�<�{�<�{�<�{�<w{�<^{�<�{�<�{�<w{�<`   `   �{�<s{�<o{�<�{�<�{�<�{�<�{�<�{�<�{�<w{�<�{�<z{�<l{�<z{�<�{�<w{�<�{�<�{�<�{�<�{�<�{�<�{�<o{�<s{�<`   `   w{�<|{�<q{�<p{�<�{�<�{�<�{�<�{�<v{�<_{�<�{�<�{�<�{�<�{�<�{�<_{�<v{�<�{�<�{�<�{�<�{�<p{�<q{�<|{�<`   `   d{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<d{�<�{�<�{�<r{�<�{�<r{�<�{�<�{�<d{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<`   `   �{�<�{�<�{�<�{�<x{�<�{�<�{�<�{�<u{�<�{�<{{�<R{�<�{�<R{�<{{�<�{�<u{�<�{�<�{�<�{�<x{�<�{�<�{�<�{�<`   `   �{�<y{�<M{�<�{�<�{�<u{�<�{�<�{�<�{�<�{�<Z{�<�{�<�{�<�{�<Z{�<�{�<�{�<�{�<�{�<u{�<�{�<�{�<M{�<y{�<`   `   �{�<�{�<b{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<y{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<b{�<�{�<`   `   �{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<f{�<f{�<�{�<e{�<H{�<e{�<�{�<f{�<f{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<`   `   �{�<�{�<�{�<�{�<n{�<�{�<k{�<�{�<�{�<j{�<�{�<�{�<�{�<�{�<�{�<j{�<�{�<�{�<k{�<�{�<n{�<�{�<�{�<�{�<`   `   w{�<g{�<�{�<~{�<w{�<�{�<i{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<i{�<�{�<w{�<~{�<�{�<g{�<`   `   {{�<�{�<�{�<�{�<v{�<�{�<v{�<p{�<�{�<�{�<�{�<Z{�<k{�<Z{�<�{�<�{�<�{�<p{�<v{�<�{�<v{�<�{�<�{�<�{�<`   `   �{�<�{�<�{�<�{�<�{�<}{�<k{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<k{�<}{�<�{�<�{�<�{�<�{�<`   `   �{�<p{�<^{�<�{�<�{�<n{�<z{�<�{�<�{�<r{�<�{�<�{�<�{�<�{�<�{�<r{�<�{�<�{�<z{�<n{�<�{�<�{�<^{�<p{�<`   `   �{�<�{�<|{�<�{�<�{�<�{�<�{�<�{�<�{�<t{�<�{�<�{�<�{�<�{�<�{�<t{�<�{�<�{�<�{�<�{�<�{�<�{�<|{�<�{�<`   `   �{�<�{�<�{�<�{�<x{�<�{�<�{�<h{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<h{�<�{�<�{�<x{�<�{�<�{�<�{�<`   `   9{�<�{�<z{�<R{�<|{�<�{�<q{�<K{�<�{�<x{�<�{�<q{�<R{�<q{�<�{�<x{�<�{�<K{�<q{�<�{�<|{�<R{�<z{�<�{�<`   `   s{�<�{�<x{�<N{�<�{�<�{�<�{�<�{�<�{�<z{�<�{�<�{�<�{�<�{�<�{�<z{�<�{�<�{�<�{�<�{�<�{�<N{�<x{�<�{�<`   `   �{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<g{�<k{�<�{�<�{�<�{�<k{�<g{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<`   `   l{�<v{�<{{�<�{�<�{�<S{�<�{�<�{�<Z{�<q{�<n{�<�{�<�{�<�{�<n{�<q{�<Z{�<�{�<�{�<S{�<�{�<�{�<{{�<v{�<`   `   �{�<{{�<m{�<�{�<k{�<7{�<�{�<�{�<d{�<�{�<�{�<{{�<�{�<{{�<�{�<�{�<d{�<�{�<�{�<7{�<k{�<�{�<m{�<{{�<`   `   �{�<�{�<r{�<�{�<�{�<�{�<�{�<�{�<e{�<q{�<h{�<�{�<�{�<�{�<h{�<q{�<e{�<�{�<�{�<�{�<�{�<�{�<r{�<�{�<`   `   n{�<u{�<�{�<�{�<�{�<�{�<�{�<p{�<j{�<a{�<~{�<�{�<�{�<�{�<~{�<a{�<j{�<p{�<�{�<�{�<�{�<�{�<�{�<u{�<`   `   �{�<�{�<�{�<�{�<w{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<w{�<�{�<�{�<�{�<`   `   �{�<�{�<�{�<~{�<�{�<�{�<�{�<�{�<�{�<�{�<x{�<s{�<�{�<s{�<x{�<�{�<�{�<�{�<�{�<�{�<�{�<~{�<�{�<�{�<`   `   ^{�<�{�<�{�<�{�<�{�<�{�<�{�<w{�<^{�<�{�<�{�<w{�<�{�<w{�<�{�<�{�<^{�<w{�<�{�<�{�<�{�<�{�<�{�<�{�<`   `   l{�<z{�<�{�<w{�<�{�<�{�<�{�<�{�<�{�<�{�<o{�<s{�<�{�<s{�<o{�<�{�<�{�<�{�<�{�<�{�<�{�<w{�<�{�<z{�<`   `   �{�<�{�<�{�<_{�<v{�<�{�<�{�<�{�<�{�<p{�<q{�<|{�<w{�<|{�<q{�<p{�<�{�<�{�<�{�<�{�<v{�<_{�<�{�<�{�<`   `   �{�<r{�<�{�<�{�<d{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<d{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<d{�<�{�<�{�<r{�<`   `   �{�<R{�<{{�<�{�<u{�<�{�<�{�<�{�<x{�<�{�<�{�<�{�<�{�<�{�<�{�<�{�<x{�<�{�<�{�<�{�<u{�<�{�<{{�<R{�<`   `   �z�<�z�<�z�<oz�<�z�<�z�<�z�< {�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�< {�<�z�<�z�<�z�<oz�<�z�<�z�<`   `   �z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<`   `   {�<�z�<{�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<{�<�z�<`   `   �z�<tz�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<tz�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<#{�<�z�<#{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<{�<�z�<�z�<�z�<�z�<�z�<{�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   {�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<"{�<�z�<�z�<�z�<�z�<�z�<"{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<	{�<�z�<�z�<�z�<�z�<�z�<	{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�< {�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�< {�<�z�<`   `   �z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<	{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<	{�<�z�<�z�<�z�<`   `   �z�<�z�<�z�< {�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�< {�<�z�<�z�<`   `   �z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�< {�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<2{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<{�<�z�<{�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�< {�<�z�<�z�<�z�<oz�<�z�<�z�<�z�<�z�<�z�<oz�<�z�<�z�<�z�< {�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<{�<�z�<{�<�z�<{�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<tz�<�z�<tz�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<#{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<#{�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   {�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<{�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<{�<�z�<�z�<`   `   �z�<�z�<�z�<"{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<"{�<�z�<�z�<`   `   �z�<�z�<�z�<	{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<	{�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�< {�<�z�<�z�<�z�< {�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<	{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<	{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�< {�<�z�<�z�<�z�<�z�<�z�< {�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `    {�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<`   `   2{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<`   `   �z�<{�<�z�<�z�<{�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<�z�<{�<�z�<�z�<{�<`   `   �y�<z�<Fz�<Zz�<"z�<	z�<Jz�<Jz�<z�<�y�<Sz�<Mz�<�y�<Mz�<Sz�<�y�<z�<Jz�<Jz�<	z�<"z�<Zz�<Fz�<z�<`   `   %z�<�y�<�y�<!z�<z�<=z�<@z�<z�<�y�<z�<z�<9z�< z�<9z�<z�<z�<�y�<z�<@z�<=z�<z�<!z�<�y�<�y�<`   `   �z�<;z�<z�<�y�<z�<z�<+z�<z�<z�<1z�<�y�<1z�<cz�<1z�<�y�<1z�<z�<z�<+z�<z�<z�<�y�<z�<;z�<`   `   z�<3z�<Sz�<.z�<%z�<�y�<Fz�<4z�<z�<Az�<�y�<7z�<)z�<7z�<�y�<Az�<z�<4z�<Fz�<�y�<%z�<.z�<Sz�<3z�<`   `   �y�<$z�<*z�<9z�<+z�<�y�<<z�<�y�<z�<Nz�<*z�<7z�<�y�<7z�<*z�<Nz�<z�<�y�<<z�<�y�<+z�<9z�<*z�<$z�<`   `   @z�<?z�<�y�<'z�</z�<Az�<;z�<�y�<Bz�<1z�<z�< z�<#z�< z�<z�<1z�<Bz�<�y�<;z�<Az�</z�<'z�<�y�<?z�<`   `   z�<-z�<z�<Dz�<z�<)z�<z�<z�<<z�<z�<0z�<-z�<Wz�<-z�<0z�<z�<<z�<z�<z�<)z�<z�<Dz�<z�<-z�<`   `   z�<Cz�< z�<mz�<z�<
z�<z�<5z�<Fz�<z�<�z�<!z�<z�<!z�<�z�<z�<Fz�<5z�<z�<
z�<z�<mz�< z�<Cz�<`   `   *z�<0z�<z�<Sz�<�y�<z�<z�<z�<Nz�<z�<bz�<z�<�y�<z�<bz�<z�<Nz�<z�<z�<z�<�y�<Sz�<z�<0z�<`   `   (z�<z�<�y�<4z�<�y�<z�<�y�<�y�<"z�<�y�<6z�<,z�<z�<,z�<6z�<�y�<"z�<�y�<�y�<z�<�y�<4z�<�y�<z�<`   `   Hz�<z�<z�<.z�<$z�<Jz�<9z�<Jz�<'z�<z�<z�<>z�<gz�<>z�<z�<z�<'z�<Jz�<9z�<Jz�<$z�<.z�<z�<z�<`   `   dz�<	z�<,z�<z�<z�<Oz�<.z�<\z�<8z�<z�<z�<z�<<z�<z�<z�<z�<8z�<\z�<.z�<Oz�<z�<z�<,z�<	z�<`   `   iz�<z�<'z�<z�<z�<2z�<�y�<-z�< z�<z�<4z�<z�<z�<z�<4z�<z�< z�<-z�<�y�<2z�<z�<z�<'z�<z�<`   `   ,z�<z�<�y�< z�<Dz�<Cz�<?z�<Nz�< z�<�y�<Bz�<Wz�<Kz�<Wz�<Bz�<�y�< z�<Nz�<?z�<Cz�<Dz�< z�<�y�<z�<`   `   �y�<)z�<z�<�y�<)z�< z�<<z�<Dz�<z�<z�<z�<	z�< z�<	z�<z�<z�<z�<Dz�<<z�< z�<)z�<�y�<z�<)z�<`   `   $z�<Jz�<>z�<�y�<z�<"z�<z�<z�<z�<%z�<z�<�y�<z�<�y�<z�<%z�<z�<z�<z�<"z�<z�<�y�<>z�<Jz�<`   `   gz�<#z�<z�<z�<z�<Dz�<>z�<(z�<z�<�y�<,z�<Xz�<Sz�<Xz�<,z�<�y�<z�<(z�<>z�<Dz�<z�<z�<z�<#z�<`   `   Gz�<�y�<�y�<z�<	z�<z�<-z�<Dz�<Rz�<Az�<=z�<.z�<�y�<.z�<=z�<Az�<Rz�<Dz�<-z�<z�<	z�<z�<�y�<�y�<`   `   ;z�<'z�<"z�<=z�<7z�<z�< z�<z�<=z�<Nz�<>z�<%z�<�y�<%z�<>z�<Nz�<=z�<z�< z�<z�<7z�<=z�<"z�<'z�<`   `   z�<z�<z�<z�<>z�<Fz�<1z�<)z�<z�<�y�<z�<?z�<,z�<?z�<z�<�y�<z�<)z�<1z�<Fz�<>z�<z�<z�<z�<`   `   �y�<�y�<�y�<
z�<z�<)z�<0z�<2z�<0z�<�y�<z�<(z�<�y�<(z�<z�<�y�<0z�<2z�<0z�<)z�<z�<
z�<�y�<�y�<`   `   'z�<z�<0z�<9z�<z�<z�<#z�<z�<-z�<*z�<Gz�<>z�<�y�<>z�<Gz�<*z�<-z�<z�<#z�<z�<z�<9z�<0z�<z�<`   `   Jz�<5z�<z�<8z�<9z�<z�<Bz�<6z�<3z�<�y�<z�<Cz�<�y�<Cz�<z�<�y�<3z�<6z�<Bz�<z�<9z�<8z�<z�<5z�<`   `   *z�<Ez�<%z�<z�<?z�<-z�</z�<z�<)z�<z�<Ez�<\z�<�y�<\z�<Ez�<z�<)z�<z�</z�<-z�<?z�<z�<%z�<Ez�<`   `   �y�<Mz�<Sz�<�y�<z�<Jz�<Jz�<	z�<"z�<Zz�<Fz�<z�<�y�<z�<Fz�<Zz�<"z�<	z�<Jz�<Jz�<z�<�y�<Sz�<Mz�<`   `    z�<9z�<z�<z�<�y�<z�<@z�<=z�<z�<!z�<�y�<�y�<%z�<�y�<�y�<!z�<z�<=z�<@z�<z�<�y�<z�<z�<9z�<`   `   cz�<1z�<�y�<1z�<z�<z�<+z�<z�<z�<�y�<z�<;z�<�z�<;z�<z�<�y�<z�<z�<+z�<z�<z�<1z�<�y�<1z�<`   `   )z�<7z�<�y�<Az�<z�<4z�<Fz�<�y�<%z�<.z�<Sz�<3z�<z�<3z�<Sz�<.z�<%z�<�y�<Fz�<4z�<z�<Az�<�y�<7z�<`   `   �y�<7z�<*z�<Nz�<z�<�y�<<z�<�y�<+z�<9z�<*z�<$z�<�y�<$z�<*z�<9z�<+z�<�y�<<z�<�y�<z�<Nz�<*z�<7z�<`   `   #z�< z�<z�<1z�<Bz�<�y�<;z�<Az�</z�<'z�<�y�<?z�<@z�<?z�<�y�<'z�</z�<Az�<;z�<�y�<Bz�<1z�<z�< z�<`   `   Wz�<-z�<0z�<z�<<z�<z�<z�<)z�<z�<Dz�<z�<-z�<z�<-z�<z�<Dz�<z�<)z�<z�<z�<<z�<z�<0z�<-z�<`   `   z�<!z�<�z�<z�<Fz�<5z�<z�<
z�<z�<mz�< z�<Cz�<z�<Cz�< z�<mz�<z�<
z�<z�<5z�<Fz�<z�<�z�<!z�<`   `   �y�<z�<bz�<z�<Nz�<z�<z�<z�<�y�<Sz�<z�<0z�<*z�<0z�<z�<Sz�<�y�<z�<z�<z�<Nz�<z�<bz�<z�<`   `   z�<,z�<6z�<�y�<"z�<�y�<�y�<z�<�y�<4z�<�y�<z�<(z�<z�<�y�<4z�<�y�<z�<�y�<�y�<"z�<�y�<6z�<,z�<`   `   gz�<>z�<z�<z�<'z�<Jz�<9z�<Jz�<$z�<.z�<z�<z�<Hz�<z�<z�<.z�<$z�<Jz�<9z�<Jz�<'z�<z�<z�<>z�<`   `   <z�<z�<z�<z�<8z�<\z�<.z�<Oz�<z�<z�<,z�<	z�<dz�<	z�<,z�<z�<z�<Oz�<.z�<\z�<8z�<z�<z�<z�<`   `   z�<z�<4z�<z�< z�<-z�<�y�<2z�<z�<z�<'z�<z�<iz�<z�<'z�<z�<z�<2z�<�y�<-z�< z�<z�<4z�<z�<`   `   Kz�<Wz�<Bz�<�y�< z�<Nz�<?z�<Cz�<Dz�< z�<�y�<z�<,z�<z�<�y�< z�<Dz�<Cz�<?z�<Nz�< z�<�y�<Bz�<Wz�<`   `    z�<	z�<z�<z�<z�<Dz�<<z�< z�<)z�<�y�<z�<)z�<�y�<)z�<z�<�y�<)z�< z�<<z�<Dz�<z�<z�<z�<	z�<`   `   z�<�y�<z�<%z�<z�<z�<z�<"z�<z�<�y�<>z�<Jz�<$z�<Jz�<>z�<�y�<z�<"z�<z�<z�<z�<%z�<z�<�y�<`   `   Sz�<Xz�<,z�<�y�<z�<(z�<>z�<Dz�<z�<z�<z�<#z�<gz�<#z�<z�<z�<z�<Dz�<>z�<(z�<z�<�y�<,z�<Xz�<`   `   �y�<.z�<=z�<Az�<Rz�<Dz�<-z�<z�<	z�<z�<�y�<�y�<Gz�<�y�<�y�<z�<	z�<z�<-z�<Dz�<Rz�<Az�<=z�<.z�<`   `   �y�<%z�<>z�<Nz�<=z�<z�< z�<z�<7z�<=z�<"z�<'z�<;z�<'z�<"z�<=z�<7z�<z�< z�<z�<=z�<Nz�<>z�<%z�<`   `   ,z�<?z�<z�<�y�<z�<)z�<1z�<Fz�<>z�<z�<z�<z�<z�<z�<z�<z�<>z�<Fz�<1z�<)z�<z�<�y�<z�<?z�<`   `   �y�<(z�<z�<�y�<0z�<2z�<0z�<)z�<z�<
z�<�y�<�y�<�y�<�y�<�y�<
z�<z�<)z�<0z�<2z�<0z�<�y�<z�<(z�<`   `   �y�<>z�<Gz�<*z�<-z�<z�<#z�<z�<z�<9z�<0z�<z�<'z�<z�<0z�<9z�<z�<z�<#z�<z�<-z�<*z�<Gz�<>z�<`   `   �y�<Cz�<z�<�y�<3z�<6z�<Bz�<z�<9z�<8z�<z�<5z�<Jz�<5z�<z�<8z�<9z�<z�<Bz�<6z�<3z�<�y�<z�<Cz�<`   `   �y�<\z�<Ez�<z�<)z�<z�</z�<-z�<?z�<z�<%z�<Ez�<*z�<Ez�<%z�<z�<?z�<-z�</z�<z�<)z�<z�<Ez�<\z�<`   `   �y�<�y�<y�<�y�<hy�<�y�<�y�<7y�<�y�<oy�<Ty�<sy�<�y�<sy�<Ty�<oy�<�y�<7y�<�y�<�y�<hy�<�y�<y�<�y�<`   `   �y�<�y�<�y�<|y�<uy�<�y�<by�<Ry�<�y�<�y�<ky�<ny�<^y�<ny�<ky�<�y�<�y�<Ry�<by�<�y�<uy�<|y�<�y�<�y�<`   `   y�<�y�<�y�<Ny�<�y�<�y�<qy�<�y�<�y�<�y�<�y�<�y�<[y�<�y�<�y�<�y�<�y�<�y�<qy�<�y�<�y�<Ny�<�y�<�y�<`   `   (y�<�y�<�y�<fy�<�y�<wy�<�y�<{y�<Dy�<sy�<�y�<�y�<}y�<�y�<�y�<sy�<Dy�<{y�<�y�<wy�<�y�<fy�<�y�<�y�<`   `   �y�<~y�<Ny�<my�<�y�<jy�<�y�<�y�<ey�<jy�<vy�<dy�<[y�<dy�<vy�<jy�<ey�<�y�<�y�<jy�<�y�<my�<Ny�<~y�<`   `   �y�<ny�<y�<�y�<xy�<�y�<xy�<�y�<�y�<�y�<�y�<jy�<|y�<jy�<�y�<�y�<�y�<�y�<xy�<�y�<xy�<�y�<y�<ny�<`   `   dy�<}y�<�y�<sy�<Dy�<�y�<?y�<�y�<ay�<cy�<�y�<cy�<�y�<cy�<�y�<cy�<ay�<�y�<?y�<�y�<Dy�<sy�<�y�<}y�<`   `   ty�<xy�<ry�<My�<Ty�<�y�<qy�<my�<�y�<yy�<My�<(y�<�y�<(y�<My�<yy�<�y�<my�<qy�<�y�<Ty�<My�<ry�<xy�<`   `   �y�<�y�<iy�<�y�<�y�<�y�<�y�<y�<�y�<�y�<Yy�<zy�<�y�<zy�<Yy�<�y�<�y�<y�<�y�<�y�<�y�<�y�<iy�<�y�<`   `   wy�<�y�<�y�<�y�<|y�<ny�<�y�<�y�<xy�<ny�<�y�<�y�<�y�<�y�<�y�<ny�<xy�<�y�<�y�<ny�<|y�<�y�<�y�<�y�<`   `   -y�<�y�<�y�<oy�<�y�<Gy�<ay�<�y�<�y�<py�<�y�<fy�<y�<fy�<�y�<py�<�y�<�y�<ay�<Gy�<�y�<oy�<�y�<�y�<`   `   (y�<�y�<�y�<xy�<�y�<ty�<Qy�<_y�<�y�<hy�<yy�<�y�<wy�<�y�<yy�<hy�<�y�<_y�<Qy�<ty�<�y�<xy�<�y�<�y�<`   `   {y�<�y�<�y�<�y�<oy�<�y�<�y�<Ry�<�y�<�y�<�y�<�y�<sy�<�y�<�y�<�y�<�y�<Ry�<�y�<�y�<oy�<�y�<�y�<�y�<`   `   �y�<�y�<y�<�y�<dy�<Xy�<�y�<^y�<�y�<�y�<�y�<by�<Uy�<by�<�y�<�y�<�y�<^y�<�y�<Xy�<dy�<�y�<y�<�y�<`   `   ay�<�y�<�y�<�y�<�y�<ey�<�y�<Gy�<~y�<�y�<fy�<by�<�y�<by�<fy�<�y�<~y�<Gy�<�y�<ey�<�y�<�y�<�y�<�y�<`   `   ey�<y�<�y�<�y�<~y�<�y�<�y�<hy�<�y�<�y�<�y�<ty�<�y�<ty�<�y�<�y�<�y�<hy�<�y�<�y�<~y�<�y�<�y�<y�<`   `   �y�<wy�<{y�<�y�<�y�<y�<qy�<�y�<�y�<�y�<�y�<�y�<y�<�y�<�y�<�y�<�y�<�y�<qy�<y�<�y�<�y�<{y�<wy�<`   `   �y�<sy�<�y�<�y�<�y�<�y�<my�<�y�<Ry�<y�<Vy�<by�<Dy�<by�<Vy�<y�<Ry�<�y�<my�<�y�<�y�<�y�<�y�<sy�<`   `   ey�<}y�<�y�<�y�<fy�<�y�<�y�<zy�<`y�<xy�<�y�<�y�<�y�<�y�<�y�<xy�<`y�<zy�<�y�<�y�<fy�<�y�<�y�<}y�<`   `   �y�<�y�<�y�<�y�<=y�<ry�<�y�<yy�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<yy�<�y�<ry�<=y�<�y�<�y�<�y�<`   `   �y�<�y�<�y�<�y�<�y�<�y�<ty�<py�<�y�<ny�<hy�<Wy�<Ty�<Wy�<hy�<ny�<�y�<py�<ty�<�y�<�y�<�y�<�y�<�y�<`   `   �y�<{y�<�y�<~y�<�y�<�y�<sy�<ty�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<ty�<sy�<�y�<�y�<~y�<�y�<{y�<`   `   Ny�<qy�<�y�<ry�<xy�<uy�<�y�<�y�<�y�<�y�<Ty�<�y�<�y�<�y�<Ty�<�y�<�y�<�y�<�y�<uy�<xy�<ry�<�y�<qy�<`   `   ]y�<qy�<�y�<�y�<�y�<Sy�<�y�<ty�<jy�<�y�<y�<ey�<�y�<ey�<y�<�y�<jy�<ty�<�y�<Sy�<�y�<�y�<�y�<qy�<`   `   �y�<sy�<Ty�<oy�<�y�<7y�<�y�<�y�<hy�<�y�<y�<�y�<�y�<�y�<y�<�y�<hy�<�y�<�y�<7y�<�y�<oy�<Ty�<sy�<`   `   ^y�<ny�<ky�<�y�<�y�<Ry�<by�<�y�<uy�<|y�<�y�<�y�<�y�<�y�<�y�<|y�<uy�<�y�<by�<Ry�<�y�<�y�<ky�<ny�<`   `   [y�<�y�<�y�<�y�<�y�<�y�<qy�<�y�<�y�<Ny�<�y�<�y�<y�<�y�<�y�<Ny�<�y�<�y�<qy�<�y�<�y�<�y�<�y�<�y�<`   `   }y�<�y�<�y�<sy�<Dy�<{y�<�y�<wy�<�y�<fy�<�y�<�y�<(y�<�y�<�y�<fy�<�y�<wy�<�y�<{y�<Dy�<sy�<�y�<�y�<`   `   [y�<dy�<vy�<jy�<ey�<�y�<�y�<jy�<�y�<my�<Ny�<~y�<�y�<~y�<Ny�<my�<�y�<jy�<�y�<�y�<ey�<jy�<vy�<dy�<`   `   |y�<jy�<�y�<�y�<�y�<�y�<xy�<�y�<xy�<�y�<y�<ny�<�y�<ny�<y�<�y�<xy�<�y�<xy�<�y�<�y�<�y�<�y�<jy�<`   `   �y�<cy�<�y�<cy�<ay�<�y�<?y�<�y�<Dy�<sy�<�y�<}y�<dy�<}y�<�y�<sy�<Dy�<�y�<?y�<�y�<ay�<cy�<�y�<cy�<`   `   �y�<(y�<My�<yy�<�y�<my�<qy�<�y�<Ty�<My�<ry�<xy�<ty�<xy�<ry�<My�<Ty�<�y�<qy�<my�<�y�<yy�<My�<(y�<`   `   �y�<zy�<Yy�<�y�<�y�<y�<�y�<�y�<�y�<�y�<iy�<�y�<�y�<�y�<iy�<�y�<�y�<�y�<�y�<y�<�y�<�y�<Yy�<zy�<`   `   �y�<�y�<�y�<ny�<xy�<�y�<�y�<ny�<|y�<�y�<�y�<�y�<wy�<�y�<�y�<�y�<|y�<ny�<�y�<�y�<xy�<ny�<�y�<�y�<`   `   y�<fy�<�y�<py�<�y�<�y�<ay�<Gy�<�y�<oy�<�y�<�y�<-y�<�y�<�y�<oy�<�y�<Gy�<ay�<�y�<�y�<py�<�y�<fy�<`   `   wy�<�y�<yy�<hy�<�y�<_y�<Qy�<ty�<�y�<xy�<�y�<�y�<(y�<�y�<�y�<xy�<�y�<ty�<Qy�<_y�<�y�<hy�<yy�<�y�<`   `   sy�<�y�<�y�<�y�<�y�<Ry�<�y�<�y�<oy�<�y�<�y�<�y�<{y�<�y�<�y�<�y�<oy�<�y�<�y�<Ry�<�y�<�y�<�y�<�y�<`   `   Uy�<by�<�y�<�y�<�y�<^y�<�y�<Xy�<dy�<�y�<y�<�y�<�y�<�y�<y�<�y�<dy�<Xy�<�y�<^y�<�y�<�y�<�y�<by�<`   `   �y�<by�<fy�<�y�<~y�<Gy�<�y�<ey�<�y�<�y�<�y�<�y�<ay�<�y�<�y�<�y�<�y�<ey�<�y�<Gy�<~y�<�y�<fy�<by�<`   `   �y�<ty�<�y�<�y�<�y�<hy�<�y�<�y�<~y�<�y�<�y�<y�<ey�<y�<�y�<�y�<~y�<�y�<�y�<hy�<�y�<�y�<�y�<ty�<`   `   y�<�y�<�y�<�y�<�y�<�y�<qy�<y�<�y�<�y�<{y�<wy�<�y�<wy�<{y�<�y�<�y�<y�<qy�<�y�<�y�<�y�<�y�<�y�<`   `   Dy�<by�<Vy�<y�<Ry�<�y�<my�<�y�<�y�<�y�<�y�<sy�<�y�<sy�<�y�<�y�<�y�<�y�<my�<�y�<Ry�<y�<Vy�<by�<`   `   �y�<�y�<�y�<xy�<`y�<zy�<�y�<�y�<fy�<�y�<�y�<}y�<ey�<}y�<�y�<�y�<fy�<�y�<�y�<zy�<`y�<xy�<�y�<�y�<`   `   �y�<�y�<�y�<�y�<�y�<yy�<�y�<ry�<=y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<=y�<ry�<�y�<yy�<�y�<�y�<�y�<�y�<`   `   Ty�<Wy�<hy�<ny�<�y�<py�<ty�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<�y�<ty�<py�<�y�<ny�<hy�<Wy�<`   `   �y�<�y�<�y�<�y�<�y�<ty�<sy�<�y�<�y�<~y�<�y�<{y�<�y�<{y�<�y�<~y�<�y�<�y�<sy�<ty�<�y�<�y�<�y�<�y�<`   `   �y�<�y�<Ty�<�y�<�y�<�y�<�y�<uy�<xy�<ry�<�y�<qy�<Ny�<qy�<�y�<ry�<xy�<uy�<�y�<�y�<�y�<�y�<Ty�<�y�<`   `   �y�<ey�<y�<�y�<jy�<ty�<�y�<Sy�<�y�<�y�<�y�<qy�<]y�<qy�<�y�<�y�<�y�<Sy�<�y�<ty�<jy�<�y�<y�<ey�<`   `   �x�<�x�<�x�<�x�<�x�<y�<�x�<y�<�x�<�x�< y�<�x�<Hy�<�x�< y�<�x�<�x�<y�<�x�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<y�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<$y�<�x�<�x�<�x�<
y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<
y�<�x�<�x�<�x�<$y�<�x�<�x�<`   `   'y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<y�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<`   `   'y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<$y�<�x�<�x�<y�<Jy�<y�<�x�<�x�<$y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<`   `   y�<�x�<�x�<�x�<y�< y�<y�<+y�<�x�<�x�<y�<�x�<�x�<�x�<y�<�x�<�x�<+y�<y�< y�<y�<�x�<�x�<�x�<`   `   y�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<y�<
y�<�x�<�x�<�x�<
y�<y�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<y�<�x�<�x�<y�<�x�<y�<�x�<�x�<0y�<�x�<�x�<�x�<�x�<�x�<0y�<�x�<�x�<y�<�x�<y�<�x�<�x�<y�<`   `   y�<y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<y�</y�<y�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<y�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<By�<y�<�x�<�x�<�x�<�x�< y�<�x�<�x�<�x�<�x�<y�<By�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   "y�<
y�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<&y�< y�<&y�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<
y�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<y�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<y�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<y�<�x�<�x�<�x�<y�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<$y�< y�<�x�<�x�<�x�<�x�<�x�<y�<$y�<	y�<y�<4y�<y�<	y�<$y�<y�<�x�<�x�<�x�<�x�<�x�< y�<$y�<`   `   �x�<�x�<�x�<�x�<y�<y�<
y�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<
y�<y�<y�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�</y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   
y�<�x�<�x�<�x�<�x�< y�<�x�<�x�<�x�<'y�<!y�<�x�<�x�<�x�<!y�<'y�<�x�<�x�<�x�< y�<�x�<�x�<�x�<�x�<`   `   $y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<y�<y�<�x�<�x�<�x�<y�<y�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<`   `   Hy�<�x�< y�<�x�<�x�<y�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<y�<�x�<�x�< y�<�x�<`   `   y�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<`   `   �x�<�x�<�x�<�x�<�x�<
y�<�x�<�x�<�x�<$y�<�x�<�x�<�x�<�x�<�x�<$y�<�x�<�x�<�x�<
y�<�x�<�x�<�x�<�x�<`   `   y�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<'y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<`   `   Jy�<y�<�x�<�x�<$y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<'y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<$y�<�x�<�x�<y�<`   `   �x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<y�<�x�<�x�<+y�<y�< y�<y�<�x�<�x�<�x�<y�<�x�<�x�<�x�<y�< y�<y�<+y�<�x�<�x�<y�<�x�<`   `   �x�<�x�<
y�<y�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<y�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<y�<
y�<�x�<`   `   �x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<`   `   �x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<`   `   �x�<�x�<�x�<0y�<�x�<�x�<y�<�x�<y�<�x�<�x�<y�<�x�<y�<�x�<�x�<y�<�x�<y�<�x�<�x�<0y�<�x�<�x�<`   `   /y�<y�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<y�<y�<y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<y�<`   `    y�<�x�<�x�<�x�<�x�<y�<By�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<By�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<`   `    y�<&y�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<
y�<"y�<
y�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<&y�<`   `   �x�<�x�<�x�<�x�<�x�<y�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<y�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<y�<�x�<`   `   4y�<y�<	y�<$y�<y�<�x�<�x�<�x�<�x�<�x�< y�<$y�<�x�<$y�< y�<�x�<�x�<�x�<�x�<�x�<y�<$y�<	y�<y�<`   `   �x�<�x�<�x�<�x�<�x�<y�<
y�<y�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<y�<
y�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<`   `   /y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<y�<�x�<�x�<�x�<�x�<`   `   y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<`   `   �x�<�x�<!y�<'y�<�x�<�x�<�x�< y�<�x�<�x�<�x�<�x�<
y�<�x�<�x�<�x�<�x�< y�<�x�<�x�<�x�<'y�<!y�<�x�<`   `   �x�<�x�<y�<y�<�x�<�x�<�x�<y�<�x�<�x�<�x�<�x�<$y�<�x�<�x�<�x�<�x�<y�<�x�<�x�<�x�<y�<y�<�x�<`   `   [x�<rx�<ex�<Bx�<�x�<\x�<!x�<cx�<Lx�<sx�<rx�<*x�<#x�<*x�<rx�<sx�<Lx�<cx�<!x�<\x�<�x�<Bx�<ex�<rx�<`   `   �x�<�x�<Rx�<ox�<�x�<mx�<\x�<dx�<vx�<�x�<wx�<Ex�<ix�<Ex�<wx�<�x�<vx�<dx�<\x�<mx�<�x�<ox�<Rx�<�x�<`   `   �x�<_x�<(x�<xx�<Jx�<mx�<ox�<Dx�<rx�<�x�<gx�<]x�<�x�<]x�<gx�<�x�<rx�<Dx�<ox�<mx�<Jx�<xx�<(x�<_x�<`   `   _x�<8x�<Gx�<~x�<7x�<sx�<dx�<Px�<�x�<�x�<yx�<Hx�<dx�<Hx�<yx�<�x�<�x�<Px�<dx�<sx�<7x�<~x�<Gx�<8x�<`   `   .x�<Tx�<�x�<�x�<_x�<�x�<�x�<ex�<bx�<fx�<zx�<Ox�<0x�<Ox�<zx�<fx�<bx�<ex�<�x�<�x�<_x�<�x�<�x�<Tx�<`   `   ax�<lx�<[x�<Ix�<_x�<Ex�<jx�<7x�<Sx�<nx�<Bx�<cx�<2x�<cx�<Bx�<nx�<Sx�<7x�<jx�<Ex�<_x�<Ix�<[x�<lx�<`   `   ~x�<ex�<8x�<7x�<px�<5x�<|x�<@x�<�x�<�x�<x�<�x�<Xx�<�x�<x�<�x�<�x�<@x�<|x�<5x�<px�<7x�<8x�<ex�<`   `   Zx�<Yx�<}x�<^x�<�x�<_x�<�x�<ex�<ex�<Kx�<9x�<�x�<;x�<�x�<9x�<Kx�<ex�<ex�<�x�<_x�<�x�<^x�<}x�<Yx�<`   `   �x�<dx�<�x�<Mx�<hx�<vx�<�x�<�x�<_x�<Ix�<vx�<�x�<�w�<�x�<vx�<Ix�<_x�<�x�<�x�<vx�<hx�<Mx�<�x�<dx�<`   `   �x�<Dx�<vx�<Yx�<ex�<�x�<^x�<�x�<wx�<Ix�<Vx�<�x�<_x�<�x�<Vx�<Ix�<wx�<�x�<^x�<�x�<ex�<Yx�<vx�<Dx�<`   `   ox�<%x�<�x�<�x�<Sx�<yx�<Dx�<Ux�<Wx�<+x�<<x�<�x�<�x�<�x�<<x�<+x�<Wx�<Ux�<Dx�<yx�<Sx�<�x�<�x�<%x�<`   `   �x�<Kx�<ox�<�x�<Ix�<=x�<Dx�<x�<px�<Zx�<jx�<2x�<x�<2x�<jx�<Zx�<px�<x�<Dx�<=x�<Ix�<�x�<ox�<Kx�<`   `   �x�<rx�<`x�<lx�<tx�<Ox�<*x�<lx�<]x�<px�<�x�<Ux�<_x�<Ux�<�x�<px�<]x�<lx�<*x�<Ox�<tx�<lx�<`x�<rx�<`   `   Kx�<gx�<�x�<Rx�<zx�<�x�<+x�<Cx�<Ox�<}x�<}x�<`x�<�x�<`x�<}x�<}x�<Ox�<Cx�<+x�<�x�<zx�<Rx�<�x�<gx�<`   `   Jx�<\x�<�x�<Sx�<Sx�<|x�<Gx�<mx�<�x�<�x�<�x�<@x�<7x�<@x�<�x�<�x�<�x�<mx�<Gx�<|x�<Sx�<Sx�<�x�<\x�<`   `   �x�<rx�<�x�<�x�<ex�<_x�<Zx�<fx�<ux�<yx�<gx�<^x�<Wx�<^x�<gx�<yx�<ux�<fx�<Zx�<_x�<ex�<�x�<�x�<rx�<`   `   ex�<ex�<qx�<~x�<sx�<x�<�x�<Ox�<Ex�<^x�<3x�<Yx�<~x�<Yx�<3x�<^x�<Ex�<Ox�<�x�<x�<sx�<~x�<qx�<ex�<`   `   [x�<Ox�<Yx�<px�<Ux�<Wx�<�x�<fx�<dx�<vx�<Yx�<mx�<zx�<mx�<Yx�<vx�<dx�<fx�<�x�<Wx�<Ux�<px�<Yx�<Ox�<`   `   �x�<hx�<rx�<�x�<px�<1x�<?x�<px�<kx�<2x�<Sx�<`x�<,x�<`x�<Sx�<2x�<kx�<px�<?x�<1x�<px�<�x�<rx�<hx�<`   `   �x�<�x�<vx�<xx�<mx�<ox�<ex�<ax�<[x�<,x�<ox�<{x�<-x�<{x�<ox�<,x�<[x�<ax�<ex�<ox�<mx�<xx�<vx�<�x�<`   `   Ux�<{x�<dx�<;x�<8x�<mx�<�x�<gx�<yx�<�x�<�x�<�x�<mx�<�x�<�x�<�x�<yx�<gx�<�x�<mx�<8x�<;x�<dx�<{x�<`   `   Cx�<ix�<rx�<�x�<gx�<Fx�<ox�<ox�<tx�<\x�<Jx�<:x�<;x�<:x�<Jx�<\x�<tx�<ox�<ox�<Fx�<gx�<�x�<rx�<ix�<`   `   mx�<ex�<ix�<�x�<}x�<kx�<^x�<ix�<Qx�<)x�<_x�<gx�<vx�<gx�<_x�<)x�<Qx�<ix�<^x�<kx�<}x�<�x�<ix�<ex�<`   `   Yx�<Kx�<Vx�<Lx�<9x�<zx�<Ex�<hx�<mx�<1x�<�x�<�x�<�x�<�x�<�x�<1x�<mx�<hx�<Ex�<zx�<9x�<Lx�<Vx�<Kx�<`   `   #x�<*x�<rx�<sx�<Lx�<cx�<!x�<\x�<�x�<Bx�<ex�<rx�<[x�<rx�<ex�<Bx�<�x�<\x�<!x�<cx�<Lx�<sx�<rx�<*x�<`   `   ix�<Ex�<wx�<�x�<vx�<dx�<\x�<mx�<�x�<ox�<Rx�<�x�<�x�<�x�<Rx�<ox�<�x�<mx�<\x�<dx�<vx�<�x�<wx�<Ex�<`   `   �x�<]x�<gx�<�x�<rx�<Dx�<ox�<mx�<Jx�<xx�<(x�<_x�<�x�<_x�<(x�<xx�<Jx�<mx�<ox�<Dx�<rx�<�x�<gx�<]x�<`   `   dx�<Hx�<yx�<�x�<�x�<Px�<dx�<sx�<7x�<~x�<Gx�<8x�<_x�<8x�<Gx�<~x�<7x�<sx�<dx�<Px�<�x�<�x�<yx�<Hx�<`   `   0x�<Ox�<zx�<fx�<bx�<ex�<�x�<�x�<_x�<�x�<�x�<Tx�<.x�<Tx�<�x�<�x�<_x�<�x�<�x�<ex�<bx�<fx�<zx�<Ox�<`   `   2x�<cx�<Bx�<nx�<Sx�<7x�<jx�<Ex�<_x�<Ix�<[x�<lx�<ax�<lx�<[x�<Ix�<_x�<Ex�<jx�<7x�<Sx�<nx�<Bx�<cx�<`   `   Xx�<�x�<x�<�x�<�x�<@x�<|x�<5x�<px�<7x�<8x�<ex�<~x�<ex�<8x�<7x�<px�<5x�<|x�<@x�<�x�<�x�<x�<�x�<`   `   ;x�<�x�<9x�<Kx�<ex�<ex�<�x�<_x�<�x�<^x�<}x�<Yx�<Zx�<Yx�<}x�<^x�<�x�<_x�<�x�<ex�<ex�<Kx�<9x�<�x�<`   `   �w�<�x�<vx�<Ix�<_x�<�x�<�x�<vx�<hx�<Mx�<�x�<dx�<�x�<dx�<�x�<Mx�<hx�<vx�<�x�<�x�<_x�<Ix�<vx�<�x�<`   `   _x�<�x�<Vx�<Ix�<wx�<�x�<^x�<�x�<ex�<Yx�<vx�<Dx�<�x�<Dx�<vx�<Yx�<ex�<�x�<^x�<�x�<wx�<Ix�<Vx�<�x�<`   `   �x�<�x�<<x�<+x�<Wx�<Ux�<Dx�<yx�<Sx�<�x�<�x�<%x�<ox�<%x�<�x�<�x�<Sx�<yx�<Dx�<Ux�<Wx�<+x�<<x�<�x�<`   `   x�<2x�<jx�<Zx�<px�<x�<Dx�<=x�<Ix�<�x�<ox�<Kx�<�x�<Kx�<ox�<�x�<Ix�<=x�<Dx�<x�<px�<Zx�<jx�<2x�<`   `   _x�<Ux�<�x�<px�<]x�<lx�<*x�<Ox�<tx�<lx�<`x�<rx�<�x�<rx�<`x�<lx�<tx�<Ox�<*x�<lx�<]x�<px�<�x�<Ux�<`   `   �x�<`x�<}x�<}x�<Ox�<Cx�<+x�<�x�<zx�<Rx�<�x�<gx�<Kx�<gx�<�x�<Rx�<zx�<�x�<+x�<Cx�<Ox�<}x�<}x�<`x�<`   `   7x�<@x�<�x�<�x�<�x�<mx�<Gx�<|x�<Sx�<Sx�<�x�<\x�<Jx�<\x�<�x�<Sx�<Sx�<|x�<Gx�<mx�<�x�<�x�<�x�<@x�<`   `   Wx�<^x�<gx�<yx�<ux�<fx�<Zx�<_x�<ex�<�x�<�x�<rx�<�x�<rx�<�x�<�x�<ex�<_x�<Zx�<fx�<ux�<yx�<gx�<^x�<`   `   ~x�<Yx�<3x�<^x�<Ex�<Ox�<�x�<x�<sx�<~x�<qx�<ex�<ex�<ex�<qx�<~x�<sx�<x�<�x�<Ox�<Ex�<^x�<3x�<Yx�<`   `   zx�<mx�<Yx�<vx�<dx�<fx�<�x�<Wx�<Ux�<px�<Yx�<Ox�<[x�<Ox�<Yx�<px�<Ux�<Wx�<�x�<fx�<dx�<vx�<Yx�<mx�<`   `   ,x�<`x�<Sx�<2x�<kx�<px�<?x�<1x�<px�<�x�<rx�<hx�<�x�<hx�<rx�<�x�<px�<1x�<?x�<px�<kx�<2x�<Sx�<`x�<`   `   -x�<{x�<ox�<,x�<[x�<ax�<ex�<ox�<mx�<xx�<vx�<�x�<�x�<�x�<vx�<xx�<mx�<ox�<ex�<ax�<[x�<,x�<ox�<{x�<`   `   mx�<�x�<�x�<�x�<yx�<gx�<�x�<mx�<8x�<;x�<dx�<{x�<Ux�<{x�<dx�<;x�<8x�<mx�<�x�<gx�<yx�<�x�<�x�<�x�<`   `   ;x�<:x�<Jx�<\x�<tx�<ox�<ox�<Fx�<gx�<�x�<rx�<ix�<Cx�<ix�<rx�<�x�<gx�<Fx�<ox�<ox�<tx�<\x�<Jx�<:x�<`   `   vx�<gx�<_x�<)x�<Qx�<ix�<^x�<kx�<}x�<�x�<ix�<ex�<mx�<ex�<ix�<�x�<}x�<kx�<^x�<ix�<Qx�<)x�<_x�<gx�<`   `   �x�<�x�<�x�<1x�<mx�<hx�<Ex�<zx�<9x�<Lx�<Vx�<Kx�<Yx�<Kx�<Vx�<Lx�<9x�<zx�<Ex�<hx�<mx�<1x�<�x�<�x�<`   `   x�<�w�<�w�<x�<�w�<�w�<x�<�w�<x�<�w�<�w�<Cx�<�w�<Cx�<�w�<�w�<x�<�w�<x�<�w�<�w�<x�<�w�<�w�<`   `   �w�<�w�<x�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<x�<�w�<`   `   �w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<`   `   �w�<x�<x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<x�<x�<`   `   �w�<x�<�w�<�w�<x�<�w�<�w�<6x�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<6x�<�w�<�w�<x�<�w�<�w�<x�<`   `   �w�<x�<�w�<�w�<x�<�w�<x�<x�<�w�<x�<x�< x�< x�< x�<x�<x�<�w�<x�<x�<�w�<x�<�w�<�w�<x�<`   `   �w�<�w�<x�<x�<�w�<�w�<�w�<�w�<x�<x�<�w�< x�<�w�< x�<�w�<x�<x�<�w�<�w�<�w�<�w�<x�<x�<�w�<`   `   �w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<	x�<�w�<	x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<	x�<�w�<�w�<�w�<x�<�w�<�w�< x�<�w�<�w�<x�<�w�<�w�<�w�<	x�<�w�<�w�<�w�<�w�<`   `   x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<%x�<x�<�w�<�w�<�w�<x�<%x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<Jx�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<Jx�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   x�<�w�<�w�<�w�<�w�<�w�<*x�<x�<�w�<�w�<�w�<�w�<-x�<�w�<�w�<�w�<�w�<x�<*x�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<x�<�w�<�w�<+x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<+x�<�w�<�w�<x�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<6x�<=x�<6x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   x�<�w�<�w�<�w�<�w�<�w�<�w�<x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<x�<x�<x�<x�<x�<x�<x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�< x�<x�<x�<x�<�w�<x�<x�<x�< x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<<x�<�w�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<<x�<`   `   �w�<Cx�<�w�<�w�<x�<�w�<x�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<x�<�w�<x�<�w�<�w�<Cx�<`   `   �w�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<x�<x�<�w�<x�<x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<x�<�w�<�w�<6x�<�w�<�w�<x�<�w�<�w�<x�<�w�<x�<�w�<�w�<x�<�w�<�w�<6x�<�w�<�w�<x�<�w�<`   `    x�< x�<x�<x�<�w�<x�<x�<�w�<x�<�w�<�w�<x�<�w�<x�<�w�<�w�<x�<�w�<x�<x�<�w�<x�<x�< x�<`   `   �w�< x�<�w�<x�<x�<�w�<�w�<�w�<�w�<x�<x�<�w�<�w�<�w�<x�<x�<�w�<�w�<�w�<�w�<x�<x�<�w�< x�<`   `   �w�<	x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<	x�<`   `    x�<�w�<�w�<x�<�w�<�w�<�w�<	x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<	x�<�w�<�w�<�w�<x�<�w�<�w�<`   `   �w�<�w�<x�<%x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<%x�<x�<�w�<`   `   �w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<`   `   �w�<�w�<x�<�w�<�w�<�w�<x�<Jx�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<Jx�<x�<�w�<�w�<�w�<x�<�w�<`   `   x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<`   `   -x�<�w�<�w�<�w�<�w�<x�<*x�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<*x�<x�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<+x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<+x�<�w�<�w�<�w�<�w�<�w�<`   `   =x�<6x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<6x�<`   `   �w�<�w�<�w�<�w�<x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<x�<x�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   x�<x�<x�<x�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<x�<x�<x�<`   `   x�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<x�<x�<x�< x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�< x�<x�<x�<x�<`   `   �w�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<x�<�w�<x�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<�w�<�w�<<x�<�w�<<x�<�w�<�w�<�w�<�w�<x�<�w�<�w�<x�<�w�<�w�<`   `   �w�<�w�<�w�<qw�<xw�<�w�<�w�<lw�<�w�<�w�<^w�<�w�<Rw�<�w�<^w�<�w�<�w�<lw�<�w�<�w�<xw�<qw�<�w�<�w�<`   `   �w�<xw�<hw�<Yw�<�w�<`w�<vw�<pw�<Ow�<rw�<�w�<�w�<Kw�<�w�<�w�<rw�<Ow�<pw�<vw�<`w�<�w�<Yw�<hw�<xw�<`   `   w�<�w�<uw�<uw�<�w�<gw�<�w�<�w�<yw�<�w�<�w�<�w�<;w�<�w�<�w�<�w�<yw�<�w�<�w�<gw�<�w�<uw�<uw�<�w�<`   `   �w�<�w�<xw�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<tw�<�w�<tw�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<xw�<�w�<`   `   nw�<[w�<hw�<ww�<cw�<�w�<Qw�<Ow�<�w�<�w�<Zw�<=w�<�w�<=w�<Zw�<�w�<�w�<Ow�<Qw�<�w�<cw�<ww�<hw�<[w�<`   `   ]w�<aw�<�w�<�w�<dw�<�w�<[w�<[w�<^w�<kw�<mw�<Tw�<�w�<Tw�<mw�<kw�<^w�<[w�<[w�<�w�<dw�<�w�<�w�<aw�<`   `   �w�<jw�<tw�<�w�<rw�<�w�<�w�<�w�<Ow�<?w�<�w�<hw�<Iw�<hw�<�w�<?w�<Ow�<�w�<�w�<�w�<rw�<�w�<tw�<jw�<`   `   �w�<�w�<`w�<w�<pw�<nw�<sw�<�w�<�w�<�w�<�w�<fw�<lw�<fw�<�w�<�w�<�w�<�w�<sw�<nw�<pw�<w�<`w�<�w�<`   `   �w�<�w�<�w�<�w�<�w�<cw�<vw�<�w�<`w�<{w�<�w�<kw�<�w�<kw�<�w�<{w�<`w�<�w�<vw�<cw�<�w�<�w�<�w�<�w�<`   `    w�<uw�<hw�<�w�<�w�<pw�<�w�<�w�<8w�<[w�<`w�<<w�<�w�<<w�<`w�<[w�<8w�<�w�<�w�<pw�<�w�<�w�<hw�<uw�<`   `   �w�<�w�<Pw�<�w�<�w�<]w�<�w�<�w�<{w�<~w�<�w�<ww�<�w�<ww�<�w�<~w�<{w�<�w�<�w�<]w�<�w�<�w�<Pw�<�w�<`   `   yw�<�w�<|w�<�w�<�w�<nw�<�w�<Iw�<�w�<kw�<Mw�<�w�<�w�<�w�<Mw�<kw�<�w�<Iw�<�w�<nw�<�w�<�w�<|w�<�w�<`   `   Bw�<{w�<�w�<�w�<�w�<Qw�<iw�<Hw�<�w�<�w�<Vw�<pw�<Kw�<pw�<Vw�<�w�<�w�<Hw�<iw�<Qw�<�w�<�w�<�w�<{w�<`   `   �w�<yw�<ow�<�w�<�w�<Iw�<nw�<�w�<�w�<�w�<�w�<�w�<*w�<�w�<�w�<�w�<�w�<�w�<nw�<Iw�<�w�<�w�<ow�<yw�<`   `   �w�<�w�<ow�<pw�<�w�<�w�<yw�<yw�<~w�<vw�<�w�<�w�<Hw�<�w�<�w�<vw�<~w�<yw�<yw�<�w�<�w�<pw�<ow�<�w�<`   `   rw�<�w�<�w�<`w�<�w�<�w�<�w�<�w�<sw�<Yw�<uw�<tw�<"w�<tw�<uw�<Yw�<sw�<�w�<�w�<�w�<�w�<`w�<�w�<�w�<`   `   Iw�<�w�<�w�<qw�<�w�<ow�<w�<�w�<�w�<zw�<�w�<vw�<Nw�<vw�<�w�<zw�<�w�<�w�<w�<ow�<�w�<qw�<�w�<�w�<`   `   {w�<�w�<�w�<�w�<�w�<�w�<_w�<|w�<xw�<kw�<|w�<~w�<�w�<~w�<|w�<kw�<xw�<|w�<_w�<�w�<�w�<�w�<�w�<�w�<`   `   �w�<�w�<�w�<cw�<�w�<�w�<�w�<�w�<dw�<�w�<nw�<Ww�<�w�<Ww�<nw�<�w�<dw�<�w�<�w�<�w�<�w�<cw�<�w�<�w�<`   `   �w�<uw�<w�<�w�<�w�<Qw�<nw�<�w�<Uw�<�w�<�w�<[w�<�w�<[w�<�w�<�w�<Uw�<�w�<nw�<Qw�<�w�<�w�<w�<uw�<`   `   {w�<mw�<�w�<�w�<�w�<>w�<ow�<�w�<\w�<pw�<zw�<w�<�w�<w�<zw�<pw�<\w�<�w�<ow�<>w�<�w�<�w�<�w�<mw�<`   `   �w�<�w�<�w�<\w�<uw�<�w�<�w�<�w�<�w�<Vw�<sw�<�w�<rw�<�w�<sw�<Vw�<�w�<�w�<�w�<�w�<uw�<\w�<�w�<�w�<`   `   ow�<�w�<�w�<rw�<iw�<ww�<gw�<hw�<hw�<gw�<�w�<�w�<hw�<�w�<�w�<gw�<hw�<hw�<gw�<ww�<iw�<rw�<�w�<�w�<`   `   ,w�<_w�<{w�<�w�<�w�<aw�<hw�<uw�<_w�<�w�<�w�<w�<�w�<w�<�w�<�w�<_w�<uw�<hw�<aw�<�w�<�w�<{w�<_w�<`   `   Rw�<�w�<^w�<�w�<�w�<lw�<�w�<�w�<xw�<qw�<�w�<�w�<�w�<�w�<�w�<qw�<xw�<�w�<�w�<lw�<�w�<�w�<^w�<�w�<`   `   Kw�<�w�<�w�<rw�<Ow�<pw�<vw�<`w�<�w�<Yw�<hw�<xw�<�w�<xw�<hw�<Yw�<�w�<`w�<vw�<pw�<Ow�<rw�<�w�<�w�<`   `   ;w�<�w�<�w�<�w�<yw�<�w�<�w�<gw�<�w�<uw�<uw�<�w�<w�<�w�<uw�<uw�<�w�<gw�<�w�<�w�<yw�<�w�<�w�<�w�<`   `   �w�<tw�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<xw�<�w�<�w�<�w�<xw�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<tw�<`   `   �w�<=w�<Zw�<�w�<�w�<Ow�<Qw�<�w�<cw�<ww�<hw�<[w�<nw�<[w�<hw�<ww�<cw�<�w�<Qw�<Ow�<�w�<�w�<Zw�<=w�<`   `   �w�<Tw�<mw�<kw�<^w�<[w�<[w�<�w�<dw�<�w�<�w�<aw�<]w�<aw�<�w�<�w�<dw�<�w�<[w�<[w�<^w�<kw�<mw�<Tw�<`   `   Iw�<hw�<�w�<?w�<Ow�<�w�<�w�<�w�<rw�<�w�<tw�<jw�<�w�<jw�<tw�<�w�<rw�<�w�<�w�<�w�<Ow�<?w�<�w�<hw�<`   `   lw�<fw�<�w�<�w�<�w�<�w�<sw�<nw�<pw�<w�<`w�<�w�<�w�<�w�<`w�<w�<pw�<nw�<sw�<�w�<�w�<�w�<�w�<fw�<`   `   �w�<kw�<�w�<{w�<`w�<�w�<vw�<cw�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<�w�<cw�<vw�<�w�<`w�<{w�<�w�<kw�<`   `   �w�<<w�<`w�<[w�<8w�<�w�<�w�<pw�<�w�<�w�<hw�<uw�< w�<uw�<hw�<�w�<�w�<pw�<�w�<�w�<8w�<[w�<`w�<<w�<`   `   �w�<ww�<�w�<~w�<{w�<�w�<�w�<]w�<�w�<�w�<Pw�<�w�<�w�<�w�<Pw�<�w�<�w�<]w�<�w�<�w�<{w�<~w�<�w�<ww�<`   `   �w�<�w�<Mw�<kw�<�w�<Iw�<�w�<nw�<�w�<�w�<|w�<�w�<yw�<�w�<|w�<�w�<�w�<nw�<�w�<Iw�<�w�<kw�<Mw�<�w�<`   `   Kw�<pw�<Vw�<�w�<�w�<Hw�<iw�<Qw�<�w�<�w�<�w�<{w�<Bw�<{w�<�w�<�w�<�w�<Qw�<iw�<Hw�<�w�<�w�<Vw�<pw�<`   `   *w�<�w�<�w�<�w�<�w�<�w�<nw�<Iw�<�w�<�w�<ow�<yw�<�w�<yw�<ow�<�w�<�w�<Iw�<nw�<�w�<�w�<�w�<�w�<�w�<`   `   Hw�<�w�<�w�<vw�<~w�<yw�<yw�<�w�<�w�<pw�<ow�<�w�<�w�<�w�<ow�<pw�<�w�<�w�<yw�<yw�<~w�<vw�<�w�<�w�<`   `   "w�<tw�<uw�<Yw�<sw�<�w�<�w�<�w�<�w�<`w�<�w�<�w�<rw�<�w�<�w�<`w�<�w�<�w�<�w�<�w�<sw�<Yw�<uw�<tw�<`   `   Nw�<vw�<�w�<zw�<�w�<�w�<w�<ow�<�w�<qw�<�w�<�w�<Iw�<�w�<�w�<qw�<�w�<ow�<w�<�w�<�w�<zw�<�w�<vw�<`   `   �w�<~w�<|w�<kw�<xw�<|w�<_w�<�w�<�w�<�w�<�w�<�w�<{w�<�w�<�w�<�w�<�w�<�w�<_w�<|w�<xw�<kw�<|w�<~w�<`   `   �w�<Ww�<nw�<�w�<dw�<�w�<�w�<�w�<�w�<cw�<�w�<�w�<�w�<�w�<�w�<cw�<�w�<�w�<�w�<�w�<dw�<�w�<nw�<Ww�<`   `   �w�<[w�<�w�<�w�<Uw�<�w�<nw�<Qw�<�w�<�w�<w�<uw�<�w�<uw�<w�<�w�<�w�<Qw�<nw�<�w�<Uw�<�w�<�w�<[w�<`   `   �w�<w�<zw�<pw�<\w�<�w�<ow�<>w�<�w�<�w�<�w�<mw�<{w�<mw�<�w�<�w�<�w�<>w�<ow�<�w�<\w�<pw�<zw�<w�<`   `   rw�<�w�<sw�<Vw�<�w�<�w�<�w�<�w�<uw�<\w�<�w�<�w�<�w�<�w�<�w�<\w�<uw�<�w�<�w�<�w�<�w�<Vw�<sw�<�w�<`   `   hw�<�w�<�w�<gw�<hw�<hw�<gw�<ww�<iw�<rw�<�w�<�w�<ow�<�w�<�w�<rw�<iw�<ww�<gw�<hw�<hw�<gw�<�w�<�w�<`   `   �w�<w�<�w�<�w�<_w�<uw�<hw�<aw�<�w�<�w�<{w�<_w�<,w�<_w�<{w�<�w�<�w�<aw�<hw�<uw�<_w�<�w�<�w�<w�<`   `   �v�<w�<"w�<w�<:w�<8w�<w�<<w�<�v�<w�<w�<w�<bw�<w�<w�<w�<�v�<<w�<w�<8w�<:w�<w�<"w�<w�<`   `   #w�<w�</w�<1w�<[w�<w�<�v�<Hw�<.w�<`w�<4w�<!w�<Zw�<!w�<4w�<`w�<.w�<Hw�<�v�<w�<[w�<1w�</w�<w�<`   `   Gw�<w�<$w�</w�< w�<w�<w�<)w�<w�<w�<�v�<w�<)w�<w�<�v�<w�<w�<)w�<w�<w�< w�</w�<$w�<w�<`   `   $w�<�v�<w�<:w�<�v�<4w�<Rw�<�v�<�v�<�v�<
w�<Pw�<<w�<Pw�<
w�<�v�<�v�<�v�<Rw�<4w�<�v�<:w�<w�<�v�<`   `   7w�<w�<Aw�<`w�<
w�<Sw�<Yw�<w�<.w�<!w�<6w�</w�<w�</w�<6w�<!w�<.w�<w�<Yw�<Sw�<
w�<`w�<Aw�<w�<`   `   Nw�<Qw�<Lw�<+w�<�v�<)w�<w�<6w�<Iw�<%w�<)w�<w�<Iw�<w�<)w�<%w�<Iw�<6w�<w�<)w�<�v�<+w�<Lw�<Qw�<`   `   w�<w�<w�<w�<w�<3w�<�v�</w�<$w�<w�<6w�</w�<�w�</w�<6w�<w�<$w�</w�<�v�<3w�<w�<w�<w�<w�<`   `   �v�<
w�<w�<6w�<2w�<Gw�<�v�<
w�<+w�<w�<w�<�v�<+w�<�v�<w�<w�<+w�<
w�<�v�<Gw�<2w�<6w�<w�<
w�<`   `   �v�<Ew�<,w�<w�<�v�<8w�<w�<�v�<=w�<w�<.w�<w�<w�<w�<.w�<w�<=w�<�v�<w�<8w�<�v�<w�<,w�<Ew�<`   `   �v�<Vw�<w�<�v�<�v�<Ew�<6w�<�v�<Uw�<w�<[w�<Jw�<�v�<Jw�<[w�<w�<Uw�<�v�<6w�<Ew�<�v�<�v�<w�<Vw�<`   `   w�<,w�<�v�<8w�<*w�<w�<w�< w�<`w�<"w�<;w�<(w�<�v�<(w�<;w�<"w�<`w�< w�<w�<w�<*w�<8w�<�v�<,w�<`   `   w�<w�<w�<Dw�<w�<�v�<*w�<+w�<Aw�<7w�<(w�<+w�<*w�<+w�<(w�<7w�<Aw�<+w�<*w�<�v�<w�<Dw�<w�<w�<`   `   )w�<%w�<(w�<w�<w�<Lw�<tw�<<w�<w�< w�< w�<w�<
w�<w�< w�< w�<w�<<w�<tw�<Lw�<w�<w�<(w�<%w�<`   `   w�<w�<1w�<�v�<5w�<^w�<w�<w�<
w�<�v�<w�<*w�<w�<*w�<w�<�v�<
w�<w�<w�<^w�<5w�<�v�<1w�<w�<`   `   �v�<w�<Cw�<w�<w�<w�<�v�<w�<Qw�<w�<�v�<=w�<cw�<=w�<�v�<w�<Qw�<w�<�v�<w�<w�<w�<Cw�<w�<`   `   	w�<w�<6w�</w�<w�<!w�<;w�<w�<w�<Aw�<w�<�v�<;w�<�v�<w�<Aw�<w�<w�<;w�<!w�<w�</w�<6w�<w�<`   `   $w�<w�<�v�<>w�<w�< w�<:w�<�v�<�v�<:w�<6w�<#w�<sw�<#w�<6w�<:w�<�v�<�v�<:w�< w�<w�<>w�<�v�<w�<`   `   w�<w�<�v�<?w�<
w�<w�<w�<w�<Aw�<!w�<%w�<5w�<dw�<5w�<%w�<!w�<Aw�<w�<w�<w�<
w�<?w�<�v�<w�<`   `   �v�<w�<w�<)w�<w�<#w�<0w�<-w�<<w�<w�<w�<�v�<�v�<�v�<w�<w�<<w�<-w�<0w�<#w�<w�<)w�<w�<w�<`   `   7w�<=w�<)w�<w�<)w�<w�<w�<w�<�v�<&w�<Rw�<?w�<w�<?w�<Rw�<&w�<�v�<w�<w�<w�<)w�<w�<)w�<=w�<`   `   7w�<w�<w�<w�< w�<w�<w�<w�<w�<Ww�<Dw�<;w�<3w�<;w�<Dw�<Ww�<w�<w�<w�<w�< w�<w�<w�<w�<`   `   w�<�v�<.w�<	w�<w�<Ow�<w�<
w�<.w�<Cw�<�v�<�v�<�v�<�v�<�v�<Cw�<.w�<
w�<w�<Ow�<w�<	w�<.w�<�v�<`   `   kw�<%w�<Pw�<"w�<!w�<Ew�<�v�<w�<5w�<(w�<w�<w�<w�<w�<w�<(w�<5w�<w�<�v�<Ew�<!w�<"w�<Pw�<%w�<`   `   hw�<w�<w�<�v�<w�<3w�<w�<Jw�<4w�<
w�<#w�<"w�<w�<"w�<#w�<
w�<4w�<Jw�<w�<3w�<w�<�v�<w�<w�<`   `   bw�<w�<w�<w�<�v�<<w�<w�<8w�<:w�<w�<"w�<w�<�v�<w�<"w�<w�<:w�<8w�<w�<<w�<�v�<w�<w�<w�<`   `   Zw�<!w�<4w�<`w�<.w�<Hw�<�v�<w�<[w�<1w�</w�<w�<#w�<w�</w�<1w�<[w�<w�<�v�<Hw�<.w�<`w�<4w�<!w�<`   `   )w�<w�<�v�<w�<w�<)w�<w�<w�< w�</w�<$w�<w�<Gw�<w�<$w�</w�< w�<w�<w�<)w�<w�<w�<�v�<w�<`   `   <w�<Pw�<
w�<�v�<�v�<�v�<Rw�<4w�<�v�<:w�<w�<�v�<$w�<�v�<w�<:w�<�v�<4w�<Rw�<�v�<�v�<�v�<
w�<Pw�<`   `   w�</w�<6w�<!w�<.w�<w�<Yw�<Sw�<
w�<`w�<Aw�<w�<7w�<w�<Aw�<`w�<
w�<Sw�<Yw�<w�<.w�<!w�<6w�</w�<`   `   Iw�<w�<)w�<%w�<Iw�<6w�<w�<)w�<�v�<+w�<Lw�<Qw�<Nw�<Qw�<Lw�<+w�<�v�<)w�<w�<6w�<Iw�<%w�<)w�<w�<`   `   �w�</w�<6w�<w�<$w�</w�<�v�<3w�<w�<w�<w�<w�<w�<w�<w�<w�<w�<3w�<�v�</w�<$w�<w�<6w�</w�<`   `   +w�<�v�<w�<w�<+w�<
w�<�v�<Gw�<2w�<6w�<w�<
w�<�v�<
w�<w�<6w�<2w�<Gw�<�v�<
w�<+w�<w�<w�<�v�<`   `   w�<w�<.w�<w�<=w�<�v�<w�<8w�<�v�<w�<,w�<Ew�<�v�<Ew�<,w�<w�<�v�<8w�<w�<�v�<=w�<w�<.w�<w�<`   `   �v�<Jw�<[w�<w�<Uw�<�v�<6w�<Ew�<�v�<�v�<w�<Vw�<�v�<Vw�<w�<�v�<�v�<Ew�<6w�<�v�<Uw�<w�<[w�<Jw�<`   `   �v�<(w�<;w�<"w�<`w�< w�<w�<w�<*w�<8w�<�v�<,w�<w�<,w�<�v�<8w�<*w�<w�<w�< w�<`w�<"w�<;w�<(w�<`   `   *w�<+w�<(w�<7w�<Aw�<+w�<*w�<�v�<w�<Dw�<w�<w�<w�<w�<w�<Dw�<w�<�v�<*w�<+w�<Aw�<7w�<(w�<+w�<`   `   
w�<w�< w�< w�<w�<<w�<tw�<Lw�<w�<w�<(w�<%w�<)w�<%w�<(w�<w�<w�<Lw�<tw�<<w�<w�< w�< w�<w�<`   `   w�<*w�<w�<�v�<
w�<w�<w�<^w�<5w�<�v�<1w�<w�<w�<w�<1w�<�v�<5w�<^w�<w�<w�<
w�<�v�<w�<*w�<`   `   cw�<=w�<�v�<w�<Qw�<w�<�v�<w�<w�<w�<Cw�<w�<�v�<w�<Cw�<w�<w�<w�<�v�<w�<Qw�<w�<�v�<=w�<`   `   ;w�<�v�<w�<Aw�<w�<w�<;w�<!w�<w�</w�<6w�<w�<	w�<w�<6w�</w�<w�<!w�<;w�<w�<w�<Aw�<w�<�v�<`   `   sw�<#w�<6w�<:w�<�v�<�v�<:w�< w�<w�<>w�<�v�<w�<$w�<w�<�v�<>w�<w�< w�<:w�<�v�<�v�<:w�<6w�<#w�<`   `   dw�<5w�<%w�<!w�<Aw�<w�<w�<w�<
w�<?w�<�v�<w�<w�<w�<�v�<?w�<
w�<w�<w�<w�<Aw�<!w�<%w�<5w�<`   `   �v�<�v�<w�<w�<<w�<-w�<0w�<#w�<w�<)w�<w�<w�<�v�<w�<w�<)w�<w�<#w�<0w�<-w�<<w�<w�<w�<�v�<`   `   w�<?w�<Rw�<&w�<�v�<w�<w�<w�<)w�<w�<)w�<=w�<7w�<=w�<)w�<w�<)w�<w�<w�<w�<�v�<&w�<Rw�<?w�<`   `   3w�<;w�<Dw�<Ww�<w�<w�<w�<w�< w�<w�<w�<w�<7w�<w�<w�<w�< w�<w�<w�<w�<w�<Ww�<Dw�<;w�<`   `   �v�<�v�<�v�<Cw�<.w�<
w�<w�<Ow�<w�<	w�<.w�<�v�<w�<�v�<.w�<	w�<w�<Ow�<w�<
w�<.w�<Cw�<�v�<�v�<`   `   w�<w�<w�<(w�<5w�<w�<�v�<Ew�<!w�<"w�<Pw�<%w�<kw�<%w�<Pw�<"w�<!w�<Ew�<�v�<w�<5w�<(w�<w�<w�<`   `   w�<"w�<#w�<
w�<4w�<Jw�<w�<3w�<w�<�v�<w�<w�<hw�<w�<w�<�v�<w�<3w�<w�<Jw�<4w�<
w�<#w�<"w�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<{v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<
w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<
w�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<w�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   w�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   {v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<
w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<
w�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   w�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<w�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<w�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<xv�<�v�<�v�<�v�<�v�<lv�<�v�<�v�<|v�<�v�<sv�<�v�<|v�<�v�<�v�<lv�<�v�<�v�<�v�<�v�<xv�<�v�<`   `   �v�<tv�<Xv�<�v�<�v�<�v�<�v�<uv�<v�<Pv�<~v�<�v�<�v�<�v�<~v�<Pv�<v�<uv�<�v�<�v�<�v�<�v�<Xv�<tv�<`   `   �v�<ov�<qv�<�v�<�v�<zv�<�v�<�v�<ev�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<ev�<�v�<�v�<zv�<�v�<�v�<qv�<ov�<`   `   ov�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<jv�<\v�<�v�<\v�<jv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   xv�<�v�<�v�<rv�<�v�<�v�<�v�<zv�<|v�<�v�<Gv�<�v�<�v�<�v�<Gv�<�v�<|v�<zv�<�v�<�v�<�v�<rv�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<cv�<wv�<�v�<yv�<�v�<�v�<�v�<yv�<�v�<wv�<cv�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<zv�<�v�<Qv�<�v�<zv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<xv�<Bv�<tv�<iv�<�v�<�v�<�v�<~v�<�v�<�v�<�v�<�v�<�v�<~v�<�v�<�v�<�v�<iv�<tv�<Bv�<xv�<�v�<`   `   �v�<zv�<|v�<�v�<�v�<pv�<�v�<�v�<Vv�<�v�<�v�<�v�<iv�<�v�<�v�<�v�<Vv�<�v�<�v�<pv�<�v�<�v�<|v�<zv�<`   `   �v�<jv�<�v�<�v�<�v�<Xv�<}v�<�v�<\v�<�v�<sv�<gv�<�v�<gv�<sv�<�v�<\v�<�v�<}v�<Xv�<�v�<�v�<�v�<jv�<`   `   �v�<mv�<�v�<Mv�<Zv�<vv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<vv�<Zv�<Mv�<�v�<mv�<`   `   �v�<�v�<�v�<pv�<�v�<�v�<uv�<�v�<~v�<�v�<�v�<nv�<yv�<nv�<�v�<�v�<~v�<�v�<uv�<�v�<�v�<pv�<�v�<�v�<`   `   sv�<sv�<�v�<�v�<�v�<�v�<_v�<�v�<�v�<nv�<[v�<rv�<rv�<rv�<[v�<nv�<�v�<�v�<_v�<�v�<�v�<�v�<�v�<sv�<`   `   Qv�<~v�<}v�<�v�<�v�<~v�<�v�<|v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<|v�<�v�<~v�<�v�<�v�<}v�<~v�<`   `   �v�<�v�<zv�<�v�<�v�<�v�<�v�<av�<jv�<�v�<�v�<�v�<Wv�<�v�<�v�<�v�<jv�<av�<�v�<�v�<�v�<�v�<zv�<�v�<`   `   _v�<�v�<�v�<�v�<�v�<�v�<Xv�<�v�<�v�<Zv�<�v�<�v�<�v�<�v�<�v�<Zv�<�v�<�v�<Xv�<�v�<�v�<�v�<�v�<�v�<`   `   �u�<^v�<�v�<xv�<�v�<�v�<Cv�<�v�<�v�<zv�<�v�<�v�<�v�<�v�<�v�<zv�<�v�<�v�<Cv�<�v�<�v�<xv�<�v�<^v�<`   `   Av�<pv�<�v�<dv�<�v�<�v�<�v�<�v�<jv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<jv�<�v�<�v�<�v�<�v�<dv�<�v�<pv�<`   `   �v�<�v�<fv�<�v�<�v�<iv�<�v�<tv�<Ev�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<Ev�<tv�<�v�<iv�<�v�<�v�<fv�<�v�<`   `   �v�<�v�<pv�<�v�<�v�<]v�<v�<�v�<�v�<�v�<�v�<uv�<�v�<uv�<�v�<�v�<�v�<�v�<v�<]v�<�v�<�v�<pv�<�v�<`   `   iv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<xv�<�v�<�v�<wv�<�v�<�v�<xv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<hv�<cv�<�v�<xv�<�v�<�v�<~v�<tv�<iv�<\v�<3v�<\v�<iv�<tv�<~v�<�v�<�v�<xv�<�v�<cv�<hv�<�v�<`   `   |v�<�v�<�v�<�v�<�v�<]v�<�v�<sv�<�v�<�v�<hv�<�v�<lv�<�v�<hv�<�v�<�v�<sv�<�v�<]v�<�v�<�v�<�v�<�v�<`   `   sv�<�v�<|v�<�v�<�v�<lv�<�v�<�v�<�v�<�v�<xv�<�v�<�v�<�v�<xv�<�v�<�v�<�v�<�v�<lv�<�v�<�v�<|v�<�v�<`   `   �v�<�v�<~v�<Pv�<v�<uv�<�v�<�v�<�v�<�v�<Xv�<tv�<�v�<tv�<Xv�<�v�<�v�<�v�<�v�<uv�<v�<Pv�<~v�<�v�<`   `   �v�<�v�<�v�<�v�<ev�<�v�<�v�<zv�<�v�<�v�<qv�<ov�<�v�<ov�<qv�<�v�<�v�<zv�<�v�<�v�<ev�<�v�<�v�<�v�<`   `   �v�<\v�<jv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<ov�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<jv�<\v�<`   `   �v�<�v�<Gv�<�v�<|v�<zv�<�v�<�v�<�v�<rv�<�v�<�v�<xv�<�v�<�v�<rv�<�v�<�v�<�v�<zv�<|v�<�v�<Gv�<�v�<`   `   �v�<�v�<yv�<�v�<wv�<cv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<cv�<wv�<�v�<yv�<�v�<`   `   Qv�<�v�<zv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<zv�<�v�<`   `   �v�<�v�<�v�<~v�<�v�<�v�<�v�<iv�<tv�<Bv�<xv�<�v�<�v�<�v�<xv�<Bv�<tv�<iv�<�v�<�v�<�v�<~v�<�v�<�v�<`   `   iv�<�v�<�v�<�v�<Vv�<�v�<�v�<pv�<�v�<�v�<|v�<zv�<�v�<zv�<|v�<�v�<�v�<pv�<�v�<�v�<Vv�<�v�<�v�<�v�<`   `   �v�<gv�<sv�<�v�<\v�<�v�<}v�<Xv�<�v�<�v�<�v�<jv�<�v�<jv�<�v�<�v�<�v�<Xv�<}v�<�v�<\v�<�v�<sv�<gv�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<vv�<Zv�<Mv�<�v�<mv�<�v�<mv�<�v�<Mv�<Zv�<vv�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   yv�<nv�<�v�<�v�<~v�<�v�<uv�<�v�<�v�<pv�<�v�<�v�<�v�<�v�<�v�<pv�<�v�<�v�<uv�<�v�<~v�<�v�<�v�<nv�<`   `   rv�<rv�<[v�<nv�<�v�<�v�<_v�<�v�<�v�<�v�<�v�<sv�<sv�<sv�<�v�<�v�<�v�<�v�<_v�<�v�<�v�<nv�<[v�<rv�<`   `   �v�<�v�<�v�<�v�<�v�<|v�<�v�<~v�<�v�<�v�<}v�<~v�<Qv�<~v�<}v�<�v�<�v�<~v�<�v�<|v�<�v�<�v�<�v�<�v�<`   `   Wv�<�v�<�v�<�v�<jv�<av�<�v�<�v�<�v�<�v�<zv�<�v�<�v�<�v�<zv�<�v�<�v�<�v�<�v�<av�<jv�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<Zv�<�v�<�v�<Xv�<�v�<�v�<�v�<�v�<�v�<_v�<�v�<�v�<�v�<�v�<�v�<Xv�<�v�<�v�<Zv�<�v�<�v�<`   `   �v�<�v�<�v�<zv�<�v�<�v�<Cv�<�v�<�v�<xv�<�v�<^v�<�u�<^v�<�v�<xv�<�v�<�v�<Cv�<�v�<�v�<zv�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<jv�<�v�<�v�<�v�<�v�<dv�<�v�<pv�<Av�<pv�<�v�<dv�<�v�<�v�<�v�<�v�<jv�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<Ev�<tv�<�v�<iv�<�v�<�v�<fv�<�v�<�v�<�v�<fv�<�v�<�v�<iv�<�v�<tv�<Ev�<�v�<�v�<�v�<`   `   �v�<uv�<�v�<�v�<�v�<�v�<v�<]v�<�v�<�v�<pv�<�v�<�v�<�v�<pv�<�v�<�v�<]v�<v�<�v�<�v�<�v�<�v�<uv�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<iv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   wv�<�v�<�v�<xv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<xv�<�v�<�v�<`   `   3v�<\v�<iv�<tv�<~v�<�v�<�v�<xv�<�v�<cv�<hv�<�v�<�v�<�v�<hv�<cv�<�v�<xv�<�v�<�v�<~v�<tv�<iv�<\v�<`   `   lv�<�v�<hv�<�v�<�v�<sv�<�v�<]v�<�v�<�v�<�v�<�v�<|v�<�v�<�v�<�v�<�v�<]v�<�v�<sv�<�v�<�v�<hv�<�v�<`   `   �u�<Pv�<Nv�<v�<Zv�<xv�<zv�<Pv�<Hv�<^v�<:v�<Qv�<�v�<Qv�<:v�<^v�<Hv�<Pv�<zv�<xv�<Zv�<v�<Nv�<Pv�<`   `   7v�<cv�<nv�<[v�<3v�<3v�<?v�<mv�<�v�<pv�<Uv�<0v�<1v�<0v�<Uv�<pv�<�v�<mv�<?v�<3v�<3v�<[v�<nv�<cv�<`   `   �v�<tv�<fv�<pv�<.v�<v�<@v�<sv�<Qv�<Ev�<yv�<Uv�<:v�<Uv�<yv�<Ev�<Qv�<sv�<@v�<v�<.v�<pv�<fv�<tv�<`   `   _v�<#v�<*v�<Cv�<Nv�<ov�<hv�<Sv�<v�<1v�<Fv�<?v�<Xv�<?v�<Fv�<1v�<v�<Sv�<hv�<ov�<Nv�<Cv�<*v�<#v�<`   `   gv�<)v�<\v�<=v�<v�<Vv�<@v�<>v�<Uv�<wv�<]v�<?v�<Bv�<?v�<]v�<wv�<Uv�<>v�<@v�<Vv�<v�<=v�<\v�<)v�<`   `   �v�<9v�<hv�<hv�<v�<\v�<Ev�<ov�<�v�<nv�<v�<]v�<"v�<]v�<v�<nv�<�v�<ov�<Ev�<\v�<v�<hv�<hv�<9v�<`   `   �v�<v�<@v�<jv�<rv�<vv�<'v�<hv�<`v�<"v�<=v�<Hv�<'v�<Hv�<=v�<"v�<`v�<hv�<'v�<vv�<rv�<jv�<@v�<v�<`   `   %v�<3v�<�v�<Kv�<rv�<tv�<v�<Mv�<lv�<Zv�<:v�<Nv�<\v�<Nv�<:v�<Zv�<lv�<Mv�<v�<tv�<rv�<Kv�<�v�<3v�<`   `   ;v�<lv�<�v�<$v�<Kv�<�v�<Nv�<Ov�<av�<�v�<Lv�<Uv�<Xv�<Uv�<Lv�<�v�<av�<Ov�<Nv�<�v�<Kv�<$v�<�v�<lv�<`   `   lv�<[v�<pv�<(v�<Uv�<rv�<bv�<Gv�<+v�<Cv�<-v�<Tv�<@v�<Tv�<-v�<Cv�<+v�<Gv�<bv�<rv�<Uv�<(v�<pv�<[v�<`   `   av�<Av�<Tv�<fv�<zv�<Iv�<Jv�<Lv�<Mv�<Gv�<=v�<dv�<*v�<dv�<=v�<Gv�<Mv�<Lv�<Jv�<Iv�<zv�<fv�<Tv�<Av�<`   `   jv�<^v�<Pv�<mv�<cv�<Cv�<Yv�<6v�<Xv�<@v�<[v�<v�<"v�<v�<[v�<@v�<Xv�<6v�<Yv�<Cv�<cv�<mv�<Pv�<^v�<`   `   [v�<pv�<0v�<>v�<;v�<fv�<�v�<<v�<Nv�<#v�<Rv�<�v�<;v�<�v�<Rv�<#v�<Nv�<<v�<�v�<fv�<;v�<>v�<0v�<pv�<`   `   Cv�<�v�<Pv�<Bv�<5v�<Av�<�v�<?v�<kv�<Mv�<Mv�<vv�<hv�<vv�<Mv�<Mv�<kv�<?v�<�v�<Av�<5v�<Bv�<Pv�<�v�<`   `   "v�<ev�<Nv�<Ov�<Nv�<-v�<Bv�<<v�<sv�<Vv�<&v�<Pv�<tv�<Pv�<&v�<Vv�<sv�<<v�<Bv�<-v�<Nv�<Ov�<Nv�<ev�<`   `   v�<Iv�<;v�<Iv�<Jv�<ev�<{v�<bv�<iv�<Yv�<"v�<8v�<@v�<8v�<"v�<Yv�<iv�<bv�<{v�<ev�<Jv�<Iv�<;v�<Iv�<`   `   w�<vv�<fv�<[v�<8v�<_v�<vv�<<v�<:v�<�v�<lv�<Xv�<.v�<Xv�<lv�<�v�<:v�<<v�<vv�<_v�<8v�<[v�<fv�<vv�<`   `   �v�<9v�<Qv�<Yv�<bv�<Jv�<Sv�<Jv�<1v�<�v�<Kv�<Nv�<Lv�<Nv�<Kv�<�v�<1v�<Jv�<Sv�<Jv�<bv�<Yv�<Qv�<9v�<`   `   lv�<Lv�<_v�<Ov�<nv�<Nv�<ev�<�v�<iv�<ev�<v�<,v�<Vv�<,v�<v�<ev�<iv�<�v�<ev�<Nv�<nv�<Ov�<_v�<Lv�<`   `   dv�<gv�<wv�<Xv�<Nv�<pv�<dv�<kv�<Bv�<Ov�<_v�<Av�<\v�<Av�<_v�<Ov�<Bv�<kv�<dv�<pv�<Nv�<Xv�<wv�<gv�<`   `   .v�<;v�<Bv�<Lv�<>v�<|v�<<v�<(v�<%v�<(v�<Wv�<?v�<�v�<?v�<Wv�<(v�<%v�<(v�<<v�<|v�<>v�<Lv�<Bv�<;v�<`   `   =v�<\v�<Mv�<Yv�<Nv�<vv�<0v�<Pv�<�v�<Nv�<*v�<$v�<�v�<$v�<*v�<Nv�<�v�<Pv�<0v�<vv�<Nv�<Yv�<Mv�<\v�<`   `   v�<Mv�<hv�<mv�<Lv�<�v�<Lv�<.v�<�v�<qv�<fv�<dv�<�v�<dv�<fv�<qv�<�v�<.v�<Lv�<�v�<Lv�<mv�<hv�<Mv�<`   `   ov�<Tv�<Xv�<Xv�<v�<av�<iv�<#v�<Bv�<2v�<|v�<�v�<Sv�<�v�<|v�<2v�<Bv�<#v�<iv�<av�<v�<Xv�<Xv�<Tv�<`   `   �v�<Qv�<:v�<^v�<Hv�<Pv�<zv�<xv�<Zv�<v�<Nv�<Pv�<�u�<Pv�<Nv�<v�<Zv�<xv�<zv�<Pv�<Hv�<^v�<:v�<Qv�<`   `   1v�<0v�<Uv�<pv�<�v�<mv�<?v�<3v�<3v�<[v�<nv�<cv�<7v�<cv�<nv�<[v�<3v�<3v�<?v�<mv�<�v�<pv�<Uv�<0v�<`   `   :v�<Uv�<yv�<Ev�<Qv�<sv�<@v�<v�<.v�<pv�<fv�<tv�<�v�<tv�<fv�<pv�<.v�<v�<@v�<sv�<Qv�<Ev�<yv�<Uv�<`   `   Xv�<?v�<Fv�<1v�<v�<Sv�<hv�<ov�<Nv�<Cv�<*v�<#v�<_v�<#v�<*v�<Cv�<Nv�<ov�<hv�<Sv�<v�<1v�<Fv�<?v�<`   `   Bv�<?v�<]v�<wv�<Uv�<>v�<@v�<Vv�<v�<=v�<\v�<)v�<gv�<)v�<\v�<=v�<v�<Vv�<@v�<>v�<Uv�<wv�<]v�<?v�<`   `   "v�<]v�<v�<nv�<�v�<ov�<Ev�<\v�<v�<hv�<hv�<9v�<�v�<9v�<hv�<hv�<v�<\v�<Ev�<ov�<�v�<nv�<v�<]v�<`   `   'v�<Hv�<=v�<"v�<`v�<hv�<'v�<vv�<rv�<jv�<@v�<v�<�v�<v�<@v�<jv�<rv�<vv�<'v�<hv�<`v�<"v�<=v�<Hv�<`   `   \v�<Nv�<:v�<Zv�<lv�<Mv�<v�<tv�<rv�<Kv�<�v�<3v�<%v�<3v�<�v�<Kv�<rv�<tv�<v�<Mv�<lv�<Zv�<:v�<Nv�<`   `   Xv�<Uv�<Lv�<�v�<av�<Ov�<Nv�<�v�<Kv�<$v�<�v�<lv�<;v�<lv�<�v�<$v�<Kv�<�v�<Nv�<Ov�<av�<�v�<Lv�<Uv�<`   `   @v�<Tv�<-v�<Cv�<+v�<Gv�<bv�<rv�<Uv�<(v�<pv�<[v�<lv�<[v�<pv�<(v�<Uv�<rv�<bv�<Gv�<+v�<Cv�<-v�<Tv�<`   `   *v�<dv�<=v�<Gv�<Mv�<Lv�<Jv�<Iv�<zv�<fv�<Tv�<Av�<av�<Av�<Tv�<fv�<zv�<Iv�<Jv�<Lv�<Mv�<Gv�<=v�<dv�<`   `   "v�<v�<[v�<@v�<Xv�<6v�<Yv�<Cv�<cv�<mv�<Pv�<^v�<jv�<^v�<Pv�<mv�<cv�<Cv�<Yv�<6v�<Xv�<@v�<[v�<v�<`   `   ;v�<�v�<Rv�<#v�<Nv�<<v�<�v�<fv�<;v�<>v�<0v�<pv�<[v�<pv�<0v�<>v�<;v�<fv�<�v�<<v�<Nv�<#v�<Rv�<�v�<`   `   hv�<vv�<Mv�<Mv�<kv�<?v�<�v�<Av�<5v�<Bv�<Pv�<�v�<Cv�<�v�<Pv�<Bv�<5v�<Av�<�v�<?v�<kv�<Mv�<Mv�<vv�<`   `   tv�<Pv�<&v�<Vv�<sv�<<v�<Bv�<-v�<Nv�<Ov�<Nv�<ev�<"v�<ev�<Nv�<Ov�<Nv�<-v�<Bv�<<v�<sv�<Vv�<&v�<Pv�<`   `   @v�<8v�<"v�<Yv�<iv�<bv�<{v�<ev�<Jv�<Iv�<;v�<Iv�<v�<Iv�<;v�<Iv�<Jv�<ev�<{v�<bv�<iv�<Yv�<"v�<8v�<`   `   .v�<Xv�<lv�<�v�<:v�<<v�<vv�<_v�<8v�<[v�<fv�<vv�<w�<vv�<fv�<[v�<8v�<_v�<vv�<<v�<:v�<�v�<lv�<Xv�<`   `   Lv�<Nv�<Kv�<�v�<1v�<Jv�<Sv�<Jv�<bv�<Yv�<Qv�<9v�<�v�<9v�<Qv�<Yv�<bv�<Jv�<Sv�<Jv�<1v�<�v�<Kv�<Nv�<`   `   Vv�<,v�<v�<ev�<iv�<�v�<ev�<Nv�<nv�<Ov�<_v�<Lv�<lv�<Lv�<_v�<Ov�<nv�<Nv�<ev�<�v�<iv�<ev�<v�<,v�<`   `   \v�<Av�<_v�<Ov�<Bv�<kv�<dv�<pv�<Nv�<Xv�<wv�<gv�<dv�<gv�<wv�<Xv�<Nv�<pv�<dv�<kv�<Bv�<Ov�<_v�<Av�<`   `   �v�<?v�<Wv�<(v�<%v�<(v�<<v�<|v�<>v�<Lv�<Bv�<;v�<.v�<;v�<Bv�<Lv�<>v�<|v�<<v�<(v�<%v�<(v�<Wv�<?v�<`   `   �v�<$v�<*v�<Nv�<�v�<Pv�<0v�<vv�<Nv�<Yv�<Mv�<\v�<=v�<\v�<Mv�<Yv�<Nv�<vv�<0v�<Pv�<�v�<Nv�<*v�<$v�<`   `   �v�<dv�<fv�<qv�<�v�<.v�<Lv�<�v�<Lv�<mv�<hv�<Mv�<v�<Mv�<hv�<mv�<Lv�<�v�<Lv�<.v�<�v�<qv�<fv�<dv�<`   `   Sv�<�v�<|v�<2v�<Bv�<#v�<iv�<av�<v�<Xv�<Xv�<Tv�<ov�<Tv�<Xv�<Xv�<v�<av�<iv�<#v�<Bv�<2v�<|v�<�v�<`   `   bv�< v�<v�<7v�<0v�<v�<v�<+v�<�u�<v�<Nv�<,v�<:v�<,v�<Nv�<v�<�u�<+v�<v�<v�<0v�<7v�<v�< v�<`   `   /v�<1v�<0v�<-v�<Cv�<[v�<'v�<v�<v�<!v�<5v�<'v�<v�<'v�<5v�<!v�<v�<v�<'v�<[v�<Cv�<-v�<0v�<1v�<`   `   �u�<v�<'v�<v�<Ev�<wv�<>v�<v�<Av�<+v�<v�<+v�<9v�<+v�<v�<+v�<Av�<v�<>v�<wv�<Ev�<v�<'v�<v�<`   `   3v�<@v�<2v�<)v�<Bv�<-v�<v�<<v�<Zv�<=v�<Dv�<Zv�<Tv�<Zv�<Dv�<=v�<Zv�<<v�<v�<-v�<Bv�<)v�<2v�<@v�<`   `   5v�<7v�<Av�<]v�<ov�<-v�<�u�<@v�<5v�<v�<@v�</v�<v�</v�<@v�<v�<5v�<@v�<�u�<-v�<ov�<]v�<Av�<7v�<`   `   v�<v�<v�<v�<Av�<Dv�<)v�<@v�<v�<�u�<v�<v�<'v�<v�<v�<�u�<v�<@v�<)v�<Dv�<Av�<v�<v�<v�<`   `   >v�<Rv�<"v�<v�<v�<v�<Kv�<1v�<�u�<Cv�<Sv�<9v�<�v�<9v�<Sv�<Cv�<�u�<1v�<Kv�<v�<v�<v�<"v�<Rv�<`   `   Pv�<;v�<&v�<Wv�<v�<v�<Xv�<)v�<v�<Hv�<1v�<v�<Gv�<v�<1v�<Hv�<v�<)v�<Xv�<v�<v�<Wv�<&v�<;v�<`   `   Dv�< v�<�u�<@v�<�u�<v�<Av�<7v�<@v�<v�<-v�<4v�<(v�<4v�<-v�<v�<@v�<7v�<Av�<v�<�u�<@v�<�u�< v�<`   `   Ev�<v�<v�<8v�<v�<v�< v�<-v�<\v�<v�<Tv�<yv�<"v�<yv�<Tv�<v�<\v�<-v�< v�<v�<v�<8v�<v�<v�<`   `   v�</v�<"v�<Bv�<Jv�<6v�<:v�<+v�<Nv�<v�<
v�<*v�<�u�<*v�<
v�<v�<Nv�<+v�<:v�<6v�<Jv�<Bv�<"v�</v�<`   `   �u�<9v�<,v�<(v�<v�< v�<.v�<v�<Rv�<Gv�<v�<1v�<Fv�<1v�<v�<Gv�<Rv�<v�<.v�< v�<v�<(v�<,v�<9v�<`   `   v�<v�<v�<Av�<#v�<v�<v�<v�<;v�<^v�<Jv�<v�<-v�<v�<Jv�<^v�<;v�<v�<v�<v�<#v�<Av�<v�<v�<`   `   5v�</v�<"v�<Pv�<bv�<7v�<v�<5v�<v�<'v�<>v�<�u�<�u�<�u�<>v�<'v�<v�<5v�<v�<7v�<bv�<Pv�<"v�</v�<`   `   v�<*v�<=v�<?v�<Qv�<&v�<�u�<Lv�<v�<4v�<\v�<%v�<Rv�<%v�<\v�<4v�<v�<Lv�<�u�<&v�<Qv�<?v�<=v�<*v�<`   `    v�<�u�<%v�<6v�<-v�<*v�<8v�<<v�<v�<8v�<Lv�<Ev�<Bv�<Ev�<Lv�<8v�<v�<<v�<8v�<*v�<-v�<6v�<%v�<�u�<`   `   Av�<�u�<!v�<>v�<&v�<v�<Av�<v�<v�<v�<v�<Bv�<v�<Bv�<v�<v�<v�<v�<Av�<v�<&v�<>v�<!v�<�u�<`   `   v�<�u�<Ev�<.v�<@v�< v�<v�<$v�<7v�<v�<v�<_v�<v�<_v�<v�<v�<7v�<$v�<v�< v�<@v�<.v�<Ev�<�u�<`   `   �u�<v�<Pv�<�u�<v�<,v�<�u�<v�<Bv�<v�<6v�<sv�<v�<sv�<6v�<v�<Bv�<v�<�u�<,v�<v�<�u�<Pv�<v�<`   `   3v�<'v�<5v�<v�<v�<:v�<v�<v�<<v�<v�<Av�<Uv�<v�<Uv�<Av�<v�<<v�<v�<v�<:v�<v�<v�<5v�<'v�<`   `   Uv�<)v�<v�<\v�<#v�<*v�<Jv�<Av�<Mv�<7v�<9v�<v�<v�<v�<9v�<7v�<Mv�<Av�<Jv�<*v�<#v�<\v�<v�<)v�<`   `   dv�<Rv�<v�<;v�<�u�<�u�<5v�<Mv�<v�<"v�<Hv�<v�<7v�<v�<Hv�<"v�<v�<Mv�<5v�<�u�<�u�<;v�<v�<Rv�<`   `   +v�<'v�<v�<Iv�<-v�<v�<&v�<Ov�<	v�<v�<Lv�< v�<,v�< v�<Lv�<v�<	v�<Ov�<&v�<v�<-v�<Iv�<v�<'v�<`   `   v�<�u�<)v�<Fv�<)v�<Nv�<v�<2v�</v�<2v�<(v�<�u�<.v�<�u�<(v�<2v�</v�<2v�<v�<Nv�<)v�<Fv�<)v�<�u�<`   `   :v�<,v�<Nv�<v�<�u�<+v�<v�<v�<0v�<7v�<v�< v�<bv�< v�<v�<7v�<0v�<v�<v�<+v�<�u�<v�<Nv�<,v�<`   `   v�<'v�<5v�<!v�<v�<v�<'v�<[v�<Cv�<-v�<0v�<1v�</v�<1v�<0v�<-v�<Cv�<[v�<'v�<v�<v�<!v�<5v�<'v�<`   `   9v�<+v�<v�<+v�<Av�<v�<>v�<wv�<Ev�<v�<'v�<v�<�u�<v�<'v�<v�<Ev�<wv�<>v�<v�<Av�<+v�<v�<+v�<`   `   Tv�<Zv�<Dv�<=v�<Zv�<<v�<v�<-v�<Bv�<)v�<2v�<@v�<3v�<@v�<2v�<)v�<Bv�<-v�<v�<<v�<Zv�<=v�<Dv�<Zv�<`   `   v�</v�<@v�<v�<5v�<@v�<�u�<-v�<ov�<]v�<Av�<7v�<5v�<7v�<Av�<]v�<ov�<-v�<�u�<@v�<5v�<v�<@v�</v�<`   `   'v�<v�<v�<�u�<v�<@v�<)v�<Dv�<Av�<v�<v�<v�<v�<v�<v�<v�<Av�<Dv�<)v�<@v�<v�<�u�<v�<v�<`   `   �v�<9v�<Sv�<Cv�<�u�<1v�<Kv�<v�<v�<v�<"v�<Rv�<>v�<Rv�<"v�<v�<v�<v�<Kv�<1v�<�u�<Cv�<Sv�<9v�<`   `   Gv�<v�<1v�<Hv�<v�<)v�<Xv�<v�<v�<Wv�<&v�<;v�<Pv�<;v�<&v�<Wv�<v�<v�<Xv�<)v�<v�<Hv�<1v�<v�<`   `   (v�<4v�<-v�<v�<@v�<7v�<Av�<v�<�u�<@v�<�u�< v�<Dv�< v�<�u�<@v�<�u�<v�<Av�<7v�<@v�<v�<-v�<4v�<`   `   "v�<yv�<Tv�<v�<\v�<-v�< v�<v�<v�<8v�<v�<v�<Ev�<v�<v�<8v�<v�<v�< v�<-v�<\v�<v�<Tv�<yv�<`   `   �u�<*v�<
v�<v�<Nv�<+v�<:v�<6v�<Jv�<Bv�<"v�</v�<v�</v�<"v�<Bv�<Jv�<6v�<:v�<+v�<Nv�<v�<
v�<*v�<`   `   Fv�<1v�<v�<Gv�<Rv�<v�<.v�< v�<v�<(v�<,v�<9v�<�u�<9v�<,v�<(v�<v�< v�<.v�<v�<Rv�<Gv�<v�<1v�<`   `   -v�<v�<Jv�<^v�<;v�<v�<v�<v�<#v�<Av�<v�<v�<v�<v�<v�<Av�<#v�<v�<v�<v�<;v�<^v�<Jv�<v�<`   `   �u�<�u�<>v�<'v�<v�<5v�<v�<7v�<bv�<Pv�<"v�</v�<5v�</v�<"v�<Pv�<bv�<7v�<v�<5v�<v�<'v�<>v�<�u�<`   `   Rv�<%v�<\v�<4v�<v�<Lv�<�u�<&v�<Qv�<?v�<=v�<*v�<v�<*v�<=v�<?v�<Qv�<&v�<�u�<Lv�<v�<4v�<\v�<%v�<`   `   Bv�<Ev�<Lv�<8v�<v�<<v�<8v�<*v�<-v�<6v�<%v�<�u�< v�<�u�<%v�<6v�<-v�<*v�<8v�<<v�<v�<8v�<Lv�<Ev�<`   `   v�<Bv�<v�<v�<v�<v�<Av�<v�<&v�<>v�<!v�<�u�<Av�<�u�<!v�<>v�<&v�<v�<Av�<v�<v�<v�<v�<Bv�<`   `   v�<_v�<v�<v�<7v�<$v�<v�< v�<@v�<.v�<Ev�<�u�<v�<�u�<Ev�<.v�<@v�< v�<v�<$v�<7v�<v�<v�<_v�<`   `   v�<sv�<6v�<v�<Bv�<v�<�u�<,v�<v�<�u�<Pv�<v�<�u�<v�<Pv�<�u�<v�<,v�<�u�<v�<Bv�<v�<6v�<sv�<`   `   v�<Uv�<Av�<v�<<v�<v�<v�<:v�<v�<v�<5v�<'v�<3v�<'v�<5v�<v�<v�<:v�<v�<v�<<v�<v�<Av�<Uv�<`   `   v�<v�<9v�<7v�<Mv�<Av�<Jv�<*v�<#v�<\v�<v�<)v�<Uv�<)v�<v�<\v�<#v�<*v�<Jv�<Av�<Mv�<7v�<9v�<v�<`   `   7v�<v�<Hv�<"v�<v�<Mv�<5v�<�u�<�u�<;v�<v�<Rv�<dv�<Rv�<v�<;v�<�u�<�u�<5v�<Mv�<v�<"v�<Hv�<v�<`   `   ,v�< v�<Lv�<v�<	v�<Ov�<&v�<v�<-v�<Iv�<v�<'v�<+v�<'v�<v�<Iv�<-v�<v�<&v�<Ov�<	v�<v�<Lv�< v�<`   `   .v�<�u�<(v�<2v�</v�<2v�<v�<Nv�<)v�<Fv�<)v�<�u�<v�<�u�<)v�<Fv�<)v�<Nv�<v�<2v�</v�<2v�<(v�<�u�<`   `   cv�<v�<v�<3v�<�u�<�u�<v�<Gv�<:v�<v�<v�<v�<�u�<v�<v�<v�<:v�<Gv�<v�<�u�<�u�<3v�<v�<v�<`   `   !v�<v�<�u�<v�<�u�<�u�<$v�</v�<&v�<v�<v�<7v�<v�<7v�<v�<v�<&v�</v�<$v�<�u�<�u�<v�<�u�<v�<`   `   �u�<v�<
v�<v�<v�<�u�<v�<�u�< v�<v�<�u�<v�<
v�<v�<�u�<v�< v�<�u�<v�<�u�<v�<v�<
v�<v�<`   `   v�<-v�<v�<v�<�u�<�u�<.v�<v�<�u�<v�<�u�<�u�<�u�<�u�<�u�<v�<�u�<v�<.v�<�u�<�u�<v�<v�<-v�<`   `   v�<!v�<�u�<�u�<�u�<v�<Bv�<v�<v�<v�<v�<v�<&v�<v�<v�<v�<v�<v�<Bv�<v�<�u�<�u�<�u�<!v�<`   `   �u�<,v�<v�<�u�<v�<v�<v�<�u�</v�<&v�<�u�<�u�<9v�<�u�<�u�<&v�</v�<�u�<v�<v�<v�<�u�<v�<,v�<`   `   �u�<Lv�<(v�<v�<v�<�u�<v�<�u�<Hv�<Sv�<v�<�u�<v�<�u�<v�<Sv�<Hv�<�u�<v�<�u�<v�<v�<(v�<Lv�<`   `   �u�<#v�<�u�<v�<7v�<v�<v�<v�<v�<�u�<v�<�u�<�u�<�u�<v�<�u�<v�<v�<v�<v�<7v�<v�<�u�<#v�<`   `   v�<v�<�u�<6v�<5v�<(v�<v�<�u�<
v�<�u�<�u�<�u�<v�<�u�<�u�<�u�<
v�<�u�<v�<(v�<5v�<6v�<�u�<v�<`   `   v�<9v�<<v�<9v�<v�<v�<�u�<�u�<v�<.v�</v�<�u�<v�<�u�</v�<.v�<v�<�u�<�u�<v�<v�<9v�<<v�<9v�<`   `   �u�<+v�<v�<�u�<�u�<v�<(v�<v�<�u�<1v�<1v�<�u�<%v�<�u�<1v�<1v�<�u�<v�<(v�<v�<�u�<�u�<v�<+v�<`   `   v�<6v�<v�<�u�<v�<*v�<'v�<!v�<�u�<v�<v�<�u�<Tv�<�u�<v�<v�<�u�<!v�<'v�<*v�<v�<�u�<v�<6v�<`   `   %v�<v�<1v�<0v�<v�</v�<�u�<(v�<v�<�u�<v�<�u�<Pv�<�u�<v�<�u�<v�<(v�<�u�</v�<v�<0v�<1v�<v�<`   `   ,v�<�u�<�u�<�u�<�u�<6v�<v�<Dv�<v�<�u�<v�<v�<bv�<v�<v�<�u�<v�<Dv�<v�<6v�<�u�<�u�<�u�<�u�<`   `   Qv�<%v�<v�<�u�<�u�<:v�<v�<-v�<�u�<�u�<v�<�u�<.v�<�u�<v�<�u�<�u�<-v�<v�<:v�<�u�<�u�<v�<%v�<`   `   v�<Lv�<Hv�<�u�<v�<v�<�u�<�u�<v�<v�< v�<�u�<�u�<�u�< v�<v�<v�<�u�<�u�<v�<v�<�u�<Hv�<Lv�<`   `   �u�<)v�<v�<�u�<v�<�u�<�u�<v�<Mv�<v�<�u�<"v�<v�<"v�<�u�<v�<Mv�<v�<�u�<�u�<v�<�u�<v�<)v�<`   `   )v�<Dv�<v�<�u�<$v�<v�<Av�<8v�<0v�<+v�<v�<v�< v�<v�<v�<+v�<0v�<8v�<Av�<v�<$v�<�u�<v�<Dv�<`   `   Nv�<2v�<v�<v�<"v�<'v�<Iv�<v�<�u�<v�<v�<�u�<�u�<�u�<v�<v�<�u�<v�<Iv�<'v�<"v�<v�<v�<2v�<`   `   /v�<v�<�u�<v�<v�<�u�<v�<v�<v�<v�<�u�<�u�<v�<�u�<�u�<v�<v�<v�<v�<�u�<v�<v�<�u�<v�<`   `   �u�<v�<v�<)v�<1v�<v�<v�<v�<7v�<&v�<�u�<v�<v�<v�<�u�<&v�<7v�<v�<v�<v�<1v�<)v�<v�<v�<`   `   �u�<v�<v�<�u�<,v�<,v�<v�<�u�<�u�<v�<0v�<>v�<v�<>v�<0v�<v�<�u�<�u�<v�<,v�<,v�<�u�<v�<v�<`   `   v�<:v�<v�<�u�<&v�<v�<v�<$v�<�u�<�u�<v�<v�<v�<v�<v�<�u�<�u�<$v�<v�<v�<&v�<�u�<v�<:v�<`   `   3v�<"v�< v�<v�<5v�<v�<�u�<Kv�<4v�<(v�<v�<�u�<(v�<�u�<v�<(v�<4v�<Kv�<�u�<v�<5v�<v�< v�<"v�<`   `   �u�<v�<v�<v�<:v�<Gv�<v�<�u�<�u�<3v�<v�<v�<cv�<v�<v�<3v�<�u�<�u�<v�<Gv�<:v�<v�<v�<v�<`   `   v�<7v�<v�<v�<&v�</v�<$v�<�u�<�u�<v�<�u�<v�<!v�<v�<�u�<v�<�u�<�u�<$v�</v�<&v�<v�<v�<7v�<`   `   
v�<v�<�u�<v�< v�<�u�<v�<�u�<v�<v�<
v�<v�<�u�<v�<
v�<v�<v�<�u�<v�<�u�< v�<v�<�u�<v�<`   `   �u�<�u�<�u�<v�<�u�<v�<.v�<�u�<�u�<v�<v�<-v�<v�<-v�<v�<v�<�u�<�u�<.v�<v�<�u�<v�<�u�<�u�<`   `   &v�<v�<v�<v�<v�<v�<Bv�<v�<�u�<�u�<�u�<!v�<v�<!v�<�u�<�u�<�u�<v�<Bv�<v�<v�<v�<v�<v�<`   `   9v�<�u�<�u�<&v�</v�<�u�<v�<v�<v�<�u�<v�<,v�<�u�<,v�<v�<�u�<v�<v�<v�<�u�</v�<&v�<�u�<�u�<`   `   v�<�u�<v�<Sv�<Hv�<�u�<v�<�u�<v�<v�<(v�<Lv�<�u�<Lv�<(v�<v�<v�<�u�<v�<�u�<Hv�<Sv�<v�<�u�<`   `   �u�<�u�<v�<�u�<v�<v�<v�<v�<7v�<v�<�u�<#v�<�u�<#v�<�u�<v�<7v�<v�<v�<v�<v�<�u�<v�<�u�<`   `   v�<�u�<�u�<�u�<
v�<�u�<v�<(v�<5v�<6v�<�u�<v�<v�<v�<�u�<6v�<5v�<(v�<v�<�u�<
v�<�u�<�u�<�u�<`   `   v�<�u�</v�<.v�<v�<�u�<�u�<v�<v�<9v�<<v�<9v�<v�<9v�<<v�<9v�<v�<v�<�u�<�u�<v�<.v�</v�<�u�<`   `   %v�<�u�<1v�<1v�<�u�<v�<(v�<v�<�u�<�u�<v�<+v�<�u�<+v�<v�<�u�<�u�<v�<(v�<v�<�u�<1v�<1v�<�u�<`   `   Tv�<�u�<v�<v�<�u�<!v�<'v�<*v�<v�<�u�<v�<6v�<v�<6v�<v�<�u�<v�<*v�<'v�<!v�<�u�<v�<v�<�u�<`   `   Pv�<�u�<v�<�u�<v�<(v�<�u�</v�<v�<0v�<1v�<v�<%v�<v�<1v�<0v�<v�</v�<�u�<(v�<v�<�u�<v�<�u�<`   `   bv�<v�<v�<�u�<v�<Dv�<v�<6v�<�u�<�u�<�u�<�u�<,v�<�u�<�u�<�u�<�u�<6v�<v�<Dv�<v�<�u�<v�<v�<`   `   .v�<�u�<v�<�u�<�u�<-v�<v�<:v�<�u�<�u�<v�<%v�<Qv�<%v�<v�<�u�<�u�<:v�<v�<-v�<�u�<�u�<v�<�u�<`   `   �u�<�u�< v�<v�<v�<�u�<�u�<v�<v�<�u�<Hv�<Lv�<v�<Lv�<Hv�<�u�<v�<v�<�u�<�u�<v�<v�< v�<�u�<`   `   v�<"v�<�u�<v�<Mv�<v�<�u�<�u�<v�<�u�<v�<)v�<�u�<)v�<v�<�u�<v�<�u�<�u�<v�<Mv�<v�<�u�<"v�<`   `    v�<v�<v�<+v�<0v�<8v�<Av�<v�<$v�<�u�<v�<Dv�<)v�<Dv�<v�<�u�<$v�<v�<Av�<8v�<0v�<+v�<v�<v�<`   `   �u�<�u�<v�<v�<�u�<v�<Iv�<'v�<"v�<v�<v�<2v�<Nv�<2v�<v�<v�<"v�<'v�<Iv�<v�<�u�<v�<v�<�u�<`   `   v�<�u�<�u�<v�<v�<v�<v�<�u�<v�<v�<�u�<v�</v�<v�<�u�<v�<v�<�u�<v�<v�<v�<v�<�u�<�u�<`   `   v�<v�<�u�<&v�<7v�<v�<v�<v�<1v�<)v�<v�<v�<�u�<v�<v�<)v�<1v�<v�<v�<v�<7v�<&v�<�u�<v�<`   `   v�<>v�<0v�<v�<�u�<�u�<v�<,v�<,v�<�u�<v�<v�<�u�<v�<v�<�u�<,v�<,v�<v�<�u�<�u�<v�<0v�<>v�<`   `   v�<v�<v�<�u�<�u�<$v�<v�<v�<&v�<�u�<v�<:v�<v�<:v�<v�<�u�<&v�<v�<v�<$v�<�u�<�u�<v�<v�<`   `   (v�<�u�<v�<(v�<4v�<Kv�<�u�<v�<5v�<v�< v�<"v�<3v�<"v�< v�<v�<5v�<v�<�u�<Kv�<4v�<(v�<v�<�u�<`   `   �u�<�u�<v�<�u�<�u�<%v�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<%v�<�u�<�u�<v�<�u�<`   `   �u�<v�<�u�<�u�< v�<v�<v�<�u�<�u�<v�<v�<v�<�u�<v�<v�<v�<�u�<�u�<v�<v�< v�<�u�<�u�<v�<`   `   Hv�<.v�<v�<v�<@v�<�u�<�u�<v�<	v�<v�<$v�<#v�<v�<#v�<$v�<v�<	v�<v�<�u�<�u�<@v�<v�<v�<.v�<`   `   �u�<�u�<�u�<"v�<9v�<0v�<v�<v�<�u�<�u�<
v�<v�<�u�<v�<
v�<�u�<�u�<v�<v�<0v�<9v�<"v�<�u�<�u�<`   `   v�<�u�<�u�<v�<�u�<v�<v�<�u�<�u�<
v�<v�<v�<v�<v�<v�<
v�<�u�<�u�<v�<v�<�u�<v�<�u�<�u�<`   `   _v�<v�<�u�<'v�<�u�<�u�<�u�<�u�<v�<�u�<v�<v�<�u�<v�<v�<�u�<v�<�u�<�u�<�u�<�u�<'v�<�u�<v�<`   `   v�<�u�<�u�<#v�<v�<v�<v�<v�<�u�<�u�<�u�<	v�<�u�<	v�<�u�<�u�<�u�<v�<v�<v�<v�<#v�<�u�<�u�<`   `   �u�<v�<�u�<�u�<�u�<v�<�u�<v�<v�<�u�<'v�<<v�<v�<<v�<'v�<�u�<v�<v�<�u�<v�<�u�<�u�<�u�<v�<`   `   �u�<$v�<v�<�u�<�u�<v�<�u�<v�</v�<v�<&v�<v�<Fv�<v�<&v�<v�</v�<v�<�u�<v�<�u�<�u�<v�<$v�<`   `   �u�<�u�<v�<�u�<�u�<v�<v�<(v�<�u�<�u�<�u�<�u�<?v�<�u�<�u�<�u�<�u�<(v�<v�<v�<�u�<�u�<v�<�u�<`   `   �u�<�u�<�u�<!v�<v�<�u�<�u�< v�<�u�<�u�<�u�<�u�<:v�<�u�<�u�<�u�<�u�< v�<�u�<�u�<v�<!v�<�u�<�u�<`   `   v�<�u�<�u�<v�<$v�<�u�<�u�<v�<v�<�u�< v�<	v�<�u�<	v�< v�<�u�<v�<v�<�u�<�u�<$v�<v�<�u�<�u�<`   `   v�<�u�<v�<�u�<�u�<�u�<�u�<�u�<v�<v�<v�<�u�<�u�<�u�<v�<v�<v�<�u�<�u�<�u�<�u�<�u�<v�<�u�<`   `   	v�<�u�<'v�<-v�<�u�<�u�<�u�<�u�< v�<0v�<v�<v�<�u�<v�<v�<0v�< v�<�u�<�u�<�u�<�u�<-v�<'v�<�u�<`   `   �u�<�u�<�u�<Rv�<v�<�u�<v�<�u�<v�<v�<�u�<�u�<�u�<�u�<�u�<v�<v�<�u�<v�<�u�<v�<Rv�<�u�<�u�<`   `   �u�<�u�<�u�<%v�<!v�< v�<(v�<�u�<v�<�u�<v�<v�<�u�<v�<v�<�u�<v�<�u�<(v�< v�<!v�<%v�<�u�<�u�<`   `   �u�<v�<�u�<v�<v�<
v�<v�<�u�<�u�<�u�<+v�<v�<v�<v�<+v�<�u�<�u�<�u�<v�<
v�<v�<v�<�u�<v�<`   `   �u�<�u�<�u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<v�<�u�<'v�<�u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<v�<�u�<�u�<`   `   �u�<�u�<�u�<6v�<�u�<�u�<�u�<v�<�u�<+v�<v�<�u�<Uv�<�u�<v�<+v�<�u�<v�<�u�<�u�<�u�<6v�<�u�<�u�<`   `   �u�<�u�<	v�<�u�<�u�<�u�<�u�<-v�<�u�<
v�<v�<v�<Pv�<v�<v�<
v�<�u�<-v�<�u�<�u�<�u�<�u�<	v�<�u�<`   `   5v�<>v�<"v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<�u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<"v�<>v�<`   `   �u�<�u�<v�<�u�<v�<v�<v�<�u�<@v�<v�<�u�<�u�<�u�<�u�<�u�<v�<@v�<�u�<v�<v�<v�<�u�<v�<�u�<`   `   �u�<�u�<!v�<v�<�u�<v�<v�<�u�<7v�< v�<�u�<%v�<�u�<%v�<�u�< v�<7v�<�u�<v�<v�<�u�<v�<!v�<�u�<`   `   v�<�u�<v�<v�<�u�<�u�<v�<�u�<�u�<�u�<v�<-v�<�u�<-v�<v�<�u�<�u�<�u�<v�<�u�<�u�<v�<v�<�u�<`   `   �u�<�u�<�u�<�u�<�u�<�u�<v�<%v�<�u�<�u�<v�<�u�<�u�<�u�<v�<�u�<�u�<%v�<v�<�u�<�u�<�u�<�u�<�u�<`   `   �u�<v�<v�<v�<�u�<�u�<v�<v�< v�<�u�<�u�<v�<�u�<v�<�u�<�u�< v�<v�<v�<�u�<�u�<v�<v�<v�<`   `   v�<#v�<$v�<v�<	v�<v�<�u�<�u�<@v�<v�<v�<.v�<Hv�<.v�<v�<v�<@v�<�u�<�u�<v�<	v�<v�<$v�<#v�<`   `   �u�<v�<
v�<�u�<�u�<v�<v�<0v�<9v�<"v�<�u�<�u�<�u�<�u�<�u�<"v�<9v�<0v�<v�<v�<�u�<�u�<
v�<v�<`   `   v�<v�<v�<
v�<�u�<�u�<v�<v�<�u�<v�<�u�<�u�<v�<�u�<�u�<v�<�u�<v�<v�<�u�<�u�<
v�<v�<v�<`   `   �u�<v�<v�<�u�<v�<�u�<�u�<�u�<�u�<'v�<�u�<v�<_v�<v�<�u�<'v�<�u�<�u�<�u�<�u�<v�<�u�<v�<v�<`   `   �u�<	v�<�u�<�u�<�u�<v�<v�<v�<v�<#v�<�u�<�u�<v�<�u�<�u�<#v�<v�<v�<v�<v�<�u�<�u�<�u�<	v�<`   `   v�<<v�<'v�<�u�<v�<v�<�u�<v�<�u�<�u�<�u�<v�<�u�<v�<�u�<�u�<�u�<v�<�u�<v�<v�<�u�<'v�<<v�<`   `   Fv�<v�<&v�<v�</v�<v�<�u�<v�<�u�<�u�<v�<$v�<�u�<$v�<v�<�u�<�u�<v�<�u�<v�</v�<v�<&v�<v�<`   `   ?v�<�u�<�u�<�u�<�u�<(v�<v�<v�<�u�<�u�<v�<�u�<�u�<�u�<v�<�u�<�u�<v�<v�<(v�<�u�<�u�<�u�<�u�<`   `   :v�<�u�<�u�<�u�<�u�< v�<�u�<�u�<v�<!v�<�u�<�u�<�u�<�u�<�u�<!v�<v�<�u�<�u�< v�<�u�<�u�<�u�<�u�<`   `   �u�<	v�< v�<�u�<v�<v�<�u�<�u�<$v�<v�<�u�<�u�<v�<�u�<�u�<v�<$v�<�u�<�u�<v�<v�<�u�< v�<	v�<`   `   �u�<�u�<v�<v�<v�<�u�<�u�<�u�<�u�<�u�<v�<�u�<v�<�u�<v�<�u�<�u�<�u�<�u�<�u�<v�<v�<v�<�u�<`   `   �u�<v�<v�<0v�< v�<�u�<�u�<�u�<�u�<-v�<'v�<�u�<	v�<�u�<'v�<-v�<�u�<�u�<�u�<�u�< v�<0v�<v�<v�<`   `   �u�<�u�<�u�<v�<v�<�u�<v�<�u�<v�<Rv�<�u�<�u�<�u�<�u�<�u�<Rv�<v�<�u�<v�<�u�<v�<v�<�u�<�u�<`   `   �u�<v�<v�<�u�<v�<�u�<(v�< v�<!v�<%v�<�u�<�u�<�u�<�u�<�u�<%v�<!v�< v�<(v�<�u�<v�<�u�<v�<v�<`   `   v�<v�<+v�<�u�<�u�<�u�<v�<
v�<v�<v�<�u�<v�<�u�<v�<�u�<v�<v�<
v�<v�<�u�<�u�<�u�<+v�<v�<`   `   'v�<�u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<v�<�u�<�u�<�u�<�u�<�u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<v�<�u�<`   `   Uv�<�u�<v�<+v�<�u�<v�<�u�<�u�<�u�<6v�<�u�<�u�<�u�<�u�<�u�<6v�<�u�<�u�<�u�<v�<�u�<+v�<v�<�u�<`   `   Pv�<v�<v�<
v�<�u�<-v�<�u�<�u�<�u�<�u�<	v�<�u�<�u�<�u�<	v�<�u�<�u�<�u�<�u�<-v�<�u�<
v�<v�<v�<`   `   �u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<"v�<>v�<5v�<>v�<"v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<`   `   �u�<�u�<�u�<v�<@v�<�u�<v�<v�<v�<�u�<v�<�u�<�u�<�u�<v�<�u�<v�<v�<v�<�u�<@v�<v�<�u�<�u�<`   `   �u�<%v�<�u�< v�<7v�<�u�<v�<v�<�u�<v�<!v�<�u�<�u�<�u�<!v�<v�<�u�<v�<v�<�u�<7v�< v�<�u�<%v�<`   `   �u�<-v�<v�<�u�<�u�<�u�<v�<�u�<�u�<v�<v�<�u�<v�<�u�<v�<v�<�u�<�u�<v�<�u�<�u�<�u�<v�<-v�<`   `   (v�<v�<�u�<v�<@v�<	v�<�u�<v�<+v�<v�<v�<.v�<8v�<.v�<v�<v�<+v�<v�<�u�<	v�<@v�<v�<�u�<v�<`   `   v�<�u�<�u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<�u�<�u�<`   `   �u�<�u�<�u�<�u�<�u�<�u�<�u�<$v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<$v�<�u�<�u�<�u�<�u�<�u�<�u�<`   `   �u�<�u�<v�<�u�<�u�<v�<�u�<v�<v�<�u�<�u�<v�<+v�<v�<�u�<�u�<v�<v�<�u�<v�<�u�<�u�<v�<�u�<`   `    v�<v�<Hv�<�u�<�u�<v�<�u�<v�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<v�<�u�<v�<�u�<�u�<Hv�<v�<`   `   v�<�u�<v�<�u�<�u�<�u�<�u�<%v�<�u�<v�<!v�<v�<v�<v�<!v�<v�<�u�<%v�<�u�<�u�<�u�<�u�<v�<�u�<`   `   v�<�u�<�u�<�u�<�u�<v�<"v�<v�<�u�<v�<	v�<v�<v�<v�<	v�<v�<�u�<v�<"v�<v�<�u�<�u�<�u�<�u�<`   `   7v�<�u�<(v�<'v�<�u�<�u�<�u�<�u�<�u�<-v�<�u�<�u�<�u�<�u�<�u�<-v�<�u�<�u�<�u�<�u�<�u�<'v�<(v�<�u�<`   `   v�<�u�<v�<=v�<(v�<�u�<�u�<�u�<�u�<v�<v�<�u�<�u�<�u�<v�<v�<�u�<�u�<�u�<�u�<(v�<=v�<v�<�u�<`   `   1v�<�u�<�u�<�u�<v�<v�< v�<�u�<�u�<�u�<v�<v�<�u�<v�<v�<�u�<�u�<�u�< v�<v�<v�<�u�<�u�<�u�<`   `   iv�<+v�<$v�<v�<�u�<v�<�u�<�u�<)v�<
v�<v�<v�<�u�<v�<v�<
v�<)v�<�u�<�u�<v�<�u�<v�<$v�<+v�<`   `   �u�<�u�< v�<v�<�u�<v�<$v�<�u�<"v�<v�<�u�<'v�<�u�<'v�<�u�<v�<"v�<�u�<$v�<v�<�u�<v�< v�<�u�<`   `   �u�<�u�<�u�<�u�<�u�<v�<Jv�<�u�<�u�<�u�<�u�<4v�<v�<4v�<�u�<�u�<�u�<�u�<Jv�<v�<�u�<�u�<�u�<�u�<`   `   v�<8v�<�u�<�u�<?v�<�u�<4v�<v�<�u�<�u�<�u�<v�<�u�<v�<�u�<�u�<�u�<v�<4v�<�u�<?v�<�u�<�u�<8v�<`   `   	v�<$v�<�u�<�u�<v�<�u�<v�<v�<�u�<�u�<�u�<v�<�u�<v�<�u�<�u�<�u�<v�<v�<�u�<v�<�u�<�u�<$v�<`   `   !v�<,v�<�u�<�u�<�u�<�u�<�u�<v�<v�<�u�<v�<v�<%v�<v�<v�<�u�<v�<v�<�u�<�u�<�u�<�u�<�u�<,v�<`   `   �u�<v�<%v�<%v�<�u�<!v�<v�<v�<*v�<�u�<v�<�u�<�u�<�u�<v�<�u�<*v�<v�<v�<!v�<�u�<%v�<%v�<v�<`   `   v�<v�<�u�<v�<�u�<5v�<�u�<v�<7v�<�u�<v�<�u�<v�<�u�<v�<�u�<7v�<v�<�u�<5v�<�u�<v�<�u�<v�<`   `   2v�<)v�<v�<�u�<�u�<9v�<�u�<v�<<v�<�u�<�u�<�u�<v�<�u�<�u�<�u�<<v�<v�<�u�<9v�<�u�<�u�<v�<)v�<`   `   �u�<�u�<v�<�u�<v�<Uv�<�u�<�u�<�u�<�u�<v�<�u�<�u�<�u�<v�<�u�<�u�<�u�<�u�<Uv�<v�<�u�<v�<�u�<`   `   �u�<�u�<�u�<�u�<v�<
v�<�u�<
v�<�u�<�u�<9v�<v�<�u�<v�<9v�<�u�<�u�<
v�<�u�<
v�<v�<�u�<�u�<�u�<`   `   iv�<�u�<�u�<(v�<v�<�u�<v�<4v�<�u�<�u�<	v�<v�<	v�<v�<	v�<�u�<�u�<4v�<v�<�u�<v�<(v�<�u�<�u�<`   `   :v�<�u�<�u�<�u�<�u�<v�<v�<�u�<�u�<v�<�u�<�u�<�u�<�u�<�u�<v�<�u�<�u�<v�<v�<�u�<�u�<�u�<�u�<`   `   v�<�u�<v�<�u�<$v�<Ov�<v�<�u�<�u�<
v�<�u�<
v�<v�<
v�<�u�<
v�<�u�<�u�<v�<Ov�<$v�<�u�<v�<�u�<`   `   8v�<.v�<v�<v�<+v�<v�<�u�<	v�<@v�<v�<�u�<v�<(v�<v�<�u�<v�<@v�<	v�<�u�<v�<+v�<v�<v�<.v�<`   `   v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<�u�<�u�<v�<�u�<�u�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<`   `   �u�<�u�<�u�<�u�<�u�<$v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<$v�<�u�<�u�<�u�<�u�<`   `   +v�<v�<�u�<�u�<v�<v�<�u�<v�<�u�<�u�<v�<�u�<�u�<�u�<v�<�u�<�u�<v�<�u�<v�<v�<�u�<�u�<v�<`   `   �u�<�u�<�u�<�u�<v�<v�<�u�<v�<�u�<�u�<Hv�<v�< v�<v�<Hv�<�u�<�u�<v�<�u�<v�<v�<�u�<�u�<�u�<`   `   v�<v�<!v�<v�<�u�<%v�<�u�<�u�<�u�<�u�<v�<�u�<v�<�u�<v�<�u�<�u�<�u�<�u�<%v�<�u�<v�<!v�<v�<`   `   v�<v�<	v�<v�<�u�<v�<"v�<v�<�u�<�u�<�u�<�u�<v�<�u�<�u�<�u�<�u�<v�<"v�<v�<�u�<v�<	v�<v�<`   `   �u�<�u�<�u�<-v�<�u�<�u�<�u�<�u�<�u�<'v�<(v�<�u�<7v�<�u�<(v�<'v�<�u�<�u�<�u�<�u�<�u�<-v�<�u�<�u�<`   `   �u�<�u�<v�<v�<�u�<�u�<�u�<�u�<(v�<=v�<v�<�u�<v�<�u�<v�<=v�<(v�<�u�<�u�<�u�<�u�<v�<v�<�u�<`   `   �u�<v�<v�<�u�<�u�<�u�< v�<v�<v�<�u�<�u�<�u�<1v�<�u�<�u�<�u�<v�<v�< v�<�u�<�u�<�u�<v�<v�<`   `   �u�<v�<v�<
v�<)v�<�u�<�u�<v�<�u�<v�<$v�<+v�<iv�<+v�<$v�<v�<�u�<v�<�u�<�u�<)v�<
v�<v�<v�<`   `   �u�<'v�<�u�<v�<"v�<�u�<$v�<v�<�u�<v�< v�<�u�<�u�<�u�< v�<v�<�u�<v�<$v�<�u�<"v�<v�<�u�<'v�<`   `   v�<4v�<�u�<�u�<�u�<�u�<Jv�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<Jv�<�u�<�u�<�u�<�u�<4v�<`   `   �u�<v�<�u�<�u�<�u�<v�<4v�<�u�<?v�<�u�<�u�<8v�<v�<8v�<�u�<�u�<?v�<�u�<4v�<v�<�u�<�u�<�u�<v�<`   `   �u�<v�<�u�<�u�<�u�<v�<v�<�u�<v�<�u�<�u�<$v�<	v�<$v�<�u�<�u�<v�<�u�<v�<v�<�u�<�u�<�u�<v�<`   `   %v�<v�<v�<�u�<v�<v�<�u�<�u�<�u�<�u�<�u�<,v�<!v�<,v�<�u�<�u�<�u�<�u�<�u�<v�<v�<�u�<v�<v�<`   `   �u�<�u�<v�<�u�<*v�<v�<v�<!v�<�u�<%v�<%v�<v�<�u�<v�<%v�<%v�<�u�<!v�<v�<v�<*v�<�u�<v�<�u�<`   `   v�<�u�<v�<�u�<7v�<v�<�u�<5v�<�u�<v�<�u�<v�<v�<v�<�u�<v�<�u�<5v�<�u�<v�<7v�<�u�<v�<�u�<`   `   v�<�u�<�u�<�u�<<v�<v�<�u�<9v�<�u�<�u�<v�<)v�<2v�<)v�<v�<�u�<�u�<9v�<�u�<v�<<v�<�u�<�u�<�u�<`   `   �u�<�u�<v�<�u�<�u�<�u�<�u�<Uv�<v�<�u�<v�<�u�<�u�<�u�<v�<�u�<v�<Uv�<�u�<�u�<�u�<�u�<v�<�u�<`   `   �u�<v�<9v�<�u�<�u�<
v�<�u�<
v�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<
v�<�u�<
v�<�u�<�u�<9v�<v�<`   `   	v�<v�<	v�<�u�<�u�<4v�<v�<�u�<v�<(v�<�u�<�u�<iv�<�u�<�u�<(v�<v�<�u�<v�<4v�<�u�<�u�<	v�<v�<`   `   �u�<�u�<�u�<v�<�u�<�u�<v�<v�<�u�<�u�<�u�<�u�<:v�<�u�<�u�<�u�<�u�<v�<v�<�u�<�u�<v�<�u�<�u�<`   `   v�<
v�<�u�<
v�<�u�<�u�<v�<Ov�<$v�<�u�<v�<�u�<v�<�u�<v�<�u�<$v�<Ov�<v�<�u�<�u�<
v�<�u�<
v�<`   `   9v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<v�<v�<v�<�u�<v�<v�<v�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<`   `   v�<�u�<#v�<#v�<�u�<v�</v�<v�<�u�<v�<v�<v�<v�<v�<v�<v�<�u�<v�</v�<v�<�u�<#v�<#v�<�u�<`   `   �u�<�u�<&v�<\v�<(v�<5v�<Bv�<v�<�u�<v�< v�<�u�<�u�<�u�< v�<v�<�u�<v�<Bv�<5v�<(v�<\v�<&v�<�u�<`   `   Hv�<#v�<�u�<-v�<#v�<v�<v�<�u�<�u�<4v�<Av�<$v�<v�<$v�<Av�<4v�<�u�<�u�<v�<v�<#v�<-v�<�u�<#v�<`   `   �u�<v�<�u�<�u�</v�<v�<Cv�<!v�<�u�<v�<v�<v�<v�<v�<v�<v�<�u�<!v�<Cv�<v�</v�<�u�<�u�<v�<`   `   �u�<v�<v�<�u�<Dv�<v�<v�<v�<�u�<v�<�u�<�u�<v�<�u�<�u�<v�<�u�<v�<v�<v�<Dv�<�u�<v�<v�<`   `   v�<(v�<@v�<�u�<(v�<�u�<�u�<�u�<	v�<9v�<�u�<v�<v�<v�<�u�<9v�<	v�<�u�<�u�<�u�<(v�<�u�<@v�<(v�<`   `   v�<�u�<v�<�u�<v�<v�<%v�<*v�<v�<v�<�u�<,v�<8v�<,v�<�u�<v�<v�<*v�<%v�<v�<v�<�u�<v�<�u�<`   `   v�<v�<v�<�u�<v�<�u�<)v�<4v�<�u�<�u�<�u�<Lv�<8v�<Lv�<�u�<�u�<�u�<4v�<)v�<�u�<v�<�u�<v�<v�<`   `   �u�<v�<!v�<�u�<v�<�u�<v�<)v�<2v�<v�<v�<;v�<
v�<;v�<v�<v�<2v�<)v�<v�<�u�<v�<�u�<!v�<v�<`   `   �u�<�u�<v�<�u�<�u�<$v�<v�<�u�<v�<v�<�u�<v�<�u�<v�<�u�<v�<v�<�u�<v�<$v�<�u�<�u�<v�<�u�<`   `   �u�<�u�<v�<v�<v�<v�<v�<�u�<�u�<v�<�u�<�u�<�u�<�u�<�u�<v�<�u�<�u�<v�<v�<v�<v�<v�<�u�<`   `   7v�<v�<v�<Cv�<>v�<�u�<�u�<v�< v�<Hv�<v�<v�<;v�<v�<v�<Hv�< v�<v�<�u�<�u�<>v�<Cv�<v�<v�<`   `   �u�<�u�< v�<v�<v�<�u�<�u�<(v�<v�<:v�< v�<v�<�u�<v�< v�<:v�<v�<(v�<�u�<�u�<v�<v�< v�<�u�<`   `   �u�<�u�<*v�<�u�<v�<Hv�<v�<v�<v�< v�<)v�<v�<�u�<v�<)v�< v�<v�<v�<v�<Hv�<v�<�u�<*v�<�u�<`   `   v�<�u�<$v�<v�<*v�<Cv�<�u�<�u�<�u�<v�< v�<�u�<)v�<�u�< v�<v�<�u�<�u�<�u�<Cv�<*v�<v�<$v�<�u�<`   `   �u�<�u�<v�<v�<$v�<v�<�u�<�u�<�u�<v�<�u�<�u�<0v�<�u�<�u�<v�<�u�<�u�<�u�<v�<$v�<v�<v�<�u�<`   `   �u�<�u�<�u�<v�<v�<v�<v�<�u�<�u�<v�<Hv�</v�<+v�</v�<Hv�<v�<�u�<�u�<v�<v�<v�<v�<�u�<�u�<`   `   	v�<v�<�u�<'v�<v�<�u�<'v�<�u�<�u�<�u�<#v�<>v�<
v�<>v�<#v�<�u�<�u�<�u�<'v�<�u�<v�<'v�<�u�<v�<`   `   v�<v�<v�<'v�<�u�<�u�<v�<�u�<#v�<v�<�u�<	v�<v�<	v�<�u�<v�<#v�<�u�<v�<�u�<�u�<'v�<v�<v�<`   `   �u�<v�<!v�< v�<�u�< v�<v�<v�<2v�<?v�<�u�< v�<Wv�< v�<�u�<?v�<2v�<v�<v�< v�<�u�< v�<!v�<v�<`   `   v�<v�<Bv�<
v�<#v�<"v�<�u�<v�<�u�<�u�<�u�<�u�<6v�<�u�<�u�<�u�<�u�<v�<�u�<"v�<#v�<
v�<Bv�<v�<`   `   �u�<7v�<Bv�<�u�<v�<�u�<�u�<5v�<�u�<v�<5v�<�u�<v�<�u�<5v�<v�<�u�<5v�<�u�<�u�<v�<�u�<Bv�<7v�<`   `   �u�< v�<v�<�u�<�u�<�u�<�u�<Cv�<v�<v�<v�<�u�<v�<�u�<v�<v�<v�<Cv�<�u�<�u�<�u�<�u�<v�< v�<`   `   �u�<v�<v�<v�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<9v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<v�<v�<v�<`   `   v�<v�<v�<v�<�u�<v�</v�<v�<�u�<#v�<#v�<�u�<v�<�u�<#v�<#v�<�u�<v�</v�<v�<�u�<v�<v�<v�<`   `   �u�<�u�< v�<v�<�u�<v�<Bv�<5v�<(v�<\v�<&v�<�u�<�u�<�u�<&v�<\v�<(v�<5v�<Bv�<v�<�u�<v�< v�<�u�<`   `   v�<$v�<Av�<4v�<�u�<�u�<v�<v�<#v�<-v�<�u�<#v�<Hv�<#v�<�u�<-v�<#v�<v�<v�<�u�<�u�<4v�<Av�<$v�<`   `   v�<v�<v�<v�<�u�<!v�<Cv�<v�</v�<�u�<�u�<v�<�u�<v�<�u�<�u�</v�<v�<Cv�<!v�<�u�<v�<v�<v�<`   `   v�<�u�<�u�<v�<�u�<v�<v�<v�<Dv�<�u�<v�<v�<�u�<v�<v�<�u�<Dv�<v�<v�<v�<�u�<v�<�u�<�u�<`   `   v�<v�<�u�<9v�<	v�<�u�<�u�<�u�<(v�<�u�<@v�<(v�<v�<(v�<@v�<�u�<(v�<�u�<�u�<�u�<	v�<9v�<�u�<v�<`   `   8v�<,v�<�u�<v�<v�<*v�<%v�<v�<v�<�u�<v�<�u�<v�<�u�<v�<�u�<v�<v�<%v�<*v�<v�<v�<�u�<,v�<`   `   8v�<Lv�<�u�<�u�<�u�<4v�<)v�<�u�<v�<�u�<v�<v�<v�<v�<v�<�u�<v�<�u�<)v�<4v�<�u�<�u�<�u�<Lv�<`   `   
v�<;v�<v�<v�<2v�<)v�<v�<�u�<v�<�u�<!v�<v�<�u�<v�<!v�<�u�<v�<�u�<v�<)v�<2v�<v�<v�<;v�<`   `   �u�<v�<�u�<v�<v�<�u�<v�<$v�<�u�<�u�<v�<�u�<�u�<�u�<v�<�u�<�u�<$v�<v�<�u�<v�<v�<�u�<v�<`   `   �u�<�u�<�u�<v�<�u�<�u�<v�<v�<v�<v�<v�<�u�<�u�<�u�<v�<v�<v�<v�<v�<�u�<�u�<v�<�u�<�u�<`   `   ;v�<v�<v�<Hv�< v�<v�<�u�<�u�<>v�<Cv�<v�<v�<7v�<v�<v�<Cv�<>v�<�u�<�u�<v�< v�<Hv�<v�<v�<`   `   �u�<v�< v�<:v�<v�<(v�<�u�<�u�<v�<v�< v�<�u�<�u�<�u�< v�<v�<v�<�u�<�u�<(v�<v�<:v�< v�<v�<`   `   �u�<v�<)v�< v�<v�<v�<v�<Hv�<v�<�u�<*v�<�u�<�u�<�u�<*v�<�u�<v�<Hv�<v�<v�<v�< v�<)v�<v�<`   `   )v�<�u�< v�<v�<�u�<�u�<�u�<Cv�<*v�<v�<$v�<�u�<v�<�u�<$v�<v�<*v�<Cv�<�u�<�u�<�u�<v�< v�<�u�<`   `   0v�<�u�<�u�<v�<�u�<�u�<�u�<v�<$v�<v�<v�<�u�<�u�<�u�<v�<v�<$v�<v�<�u�<�u�<�u�<v�<�u�<�u�<`   `   +v�</v�<Hv�<v�<�u�<�u�<v�<v�<v�<v�<�u�<�u�<�u�<�u�<�u�<v�<v�<v�<v�<�u�<�u�<v�<Hv�</v�<`   `   
v�<>v�<#v�<�u�<�u�<�u�<'v�<�u�<v�<'v�<�u�<v�<	v�<v�<�u�<'v�<v�<�u�<'v�<�u�<�u�<�u�<#v�<>v�<`   `   v�<	v�<�u�<v�<#v�<�u�<v�<�u�<�u�<'v�<v�<v�<v�<v�<v�<'v�<�u�<�u�<v�<�u�<#v�<v�<�u�<	v�<`   `   Wv�< v�<�u�<?v�<2v�<v�<v�< v�<�u�< v�<!v�<v�<�u�<v�<!v�< v�<�u�< v�<v�<v�<2v�<?v�<�u�< v�<`   `   6v�<�u�<�u�<�u�<�u�<v�<�u�<"v�<#v�<
v�<Bv�<v�<v�<v�<Bv�<
v�<#v�<"v�<�u�<v�<�u�<�u�<�u�<�u�<`   `   v�<�u�<5v�<v�<�u�<5v�<�u�<�u�<v�<�u�<Bv�<7v�<�u�<7v�<Bv�<�u�<v�<�u�<�u�<5v�<�u�<v�<5v�<�u�<`   `   v�<�u�<v�<v�<v�<Cv�<�u�<�u�<�u�<�u�<v�< v�<�u�< v�<v�<�u�<�u�<�u�<�u�<Cv�<v�<v�<v�<�u�<`   `   �u�<v�<Mv�<!v�<v�<v�<Dv�<*v�<v�<4v�<v�<v�<,v�<v�<v�<4v�<v�<*v�<Dv�<v�<v�<!v�<Mv�<v�<`   `   v�<Dv�<&v�<�u�<:v�<*v�<v�<4v�<(v�<&v�<*v�<2v�<Jv�<2v�<*v�<&v�<(v�<4v�<v�<*v�<:v�<�u�<&v�<Dv�<`   `    v�<;v�<�u�<�u�<2v�< v�<�u�<"v�<Lv�<�u�<v�<&v�<>v�<&v�<v�<�u�<Lv�<"v�<�u�< v�<2v�<�u�<�u�<;v�<`   `   v�<6v�<	v�<8v�<�u�<�u�<v�<v�<Pv�<�u�<�u�<v�<�u�<v�<�u�<�u�<Pv�<v�<v�<�u�<�u�<8v�<	v�<6v�<`   `   v�<,v�<v�<Iv�<v�<�u�<Vv�<v�<Fv�<#v�<(v�<>v�<v�<>v�<(v�<#v�<Fv�<v�<Vv�<�u�<v�<Iv�<v�<,v�<`   `   :v�<<v�<v�<*v�<v�<	v�<2v�<v�<9v�<v�<v�<Ev�<!v�<Ev�<v�<v�<9v�<v�<2v�<	v�<v�<*v�<v�<<v�<`   `   =v�< v�<2v�<9v�<*v�<v�<v�<?v�<:v�<�u�<*v�<.v�<�u�<.v�<*v�<�u�<:v�<?v�<v�<v�<*v�<9v�<2v�< v�<`   `   v�<�u�<*v�<+v�<.v�<?v�<,v�< v�<v�<v�<Tv�<Iv�<�u�<Iv�<Tv�<v�<v�< v�<,v�<?v�<.v�<+v�<*v�<�u�<`   `   /v�<>v�<0v�<v�<v�<v�<v�<�u�<v�<;v�<!v�<v�<�u�<v�<!v�<;v�<v�<�u�<v�<v�<v�<v�<0v�<>v�<`   `   v�<Qv�<Bv�<Iv�<Jv�<v�<v�<v�<7v�<@v�<�u�<�u�<v�<�u�<�u�<@v�<7v�<v�<v�<v�<Jv�<Iv�<Bv�<Qv�<`   `   v�<)v�<v�<Cv�<Cv�<v�<v�<6v�<v�<v�<2v�<8v�<yv�<8v�<2v�<v�<v�<6v�<v�<v�<Cv�<Cv�<v�<)v�<`   `   fv�<6v�<�u�<v�<v�<v�<v�<av�<v�<v�<_v�<v�<Fv�<v�<_v�<v�<v�<av�<v�<v�<v�<v�<�u�<6v�<`   `   Ov�<v�<v�<v�< v�<av�<.v�<Qv�<'v�<v�<5v�<�u�<v�<�u�<5v�<v�<'v�<Qv�<.v�<av�< v�<v�<v�<v�<`   `   Gv�<�u�<#v�<v�<�u�<cv�<+v�<	v�<v�<�u�<�u�<&v�<Lv�<&v�<�u�<�u�<v�<	v�<+v�<cv�<�u�<v�<#v�<�u�<`   `   �v�<v�<@v�<>v�<�u�<-v�<v�<v�<+v�<
v�<v�<9v�<%v�<9v�<v�<
v�<+v�<v�<v�<-v�<�u�<>v�<@v�<v�<`   `   uv�<v�<v�<9v�<v�<v�<5v�<_v�<'v�<+v�<4v�<.v�<v�<.v�<4v�<+v�<'v�<_v�<5v�<v�<v�<9v�<v�<v�<`   `   av�<?v�<v�<�u�<v�<�u�<Nv�<jv�<v�<v�<v�<-v�<Tv�<-v�<v�<v�<v�<jv�<Nv�<�u�<v�<�u�<v�<?v�<`   `   5v�<uv�<^v�<v�<+v�<v�<Bv�<.v�<"v�<@v�<�u�<v�<�u�<v�<�u�<@v�<"v�<.v�<Bv�<v�<+v�<v�<^v�<uv�<`   `   �u�<v�<v�<Fv�<_v�<v�<Vv�<v�<5v�<Gv�<
v�<v�<�u�<v�<
v�<Gv�<5v�<v�<Vv�<v�<_v�<Fv�<v�<v�<`   `   6v�</v�<�u�<0v�<Gv�<v�<Wv�<%v�<v�<"v�<,v�<]v�<0v�<]v�<,v�<"v�<v�<%v�<Wv�<v�<Gv�<0v�<�u�</v�<`   `   Yv�<Rv�<v�<v�<v�<5v�<.v�<v�<v�<v�<,v�<)v�<v�<)v�<,v�<v�<v�<v�<.v�<5v�<v�<v�<v�<Rv�<`   `   �u�<�u�<�u�<�u�<v�<av�<v�<�u�<8v�<v�<)v�< v�<�u�< v�<)v�<v�<8v�<�u�<v�<av�<v�<�u�<�u�<�u�<`   `   +v�<%v�<
v�<Mv�<>v�<2v�<v�<v�<-v�<v�<;v�<Dv�<Tv�<Dv�<;v�<v�<-v�<v�<v�<2v�<>v�<Mv�<
v�<%v�<`   `   _v�<Cv�<v�<gv�<8v�<v�<Mv�<)v�<v�<"v�<<v�< v�<2v�< v�<<v�<"v�<v�<)v�<Mv�<v�<8v�<gv�<v�<Cv�<`   `   ,v�<v�<v�<4v�<v�<*v�<Dv�<v�<v�<!v�<Mv�<v�<�u�<v�<Mv�<!v�<v�<v�<Dv�<*v�<v�<4v�<v�<v�<`   `   Jv�<2v�<*v�<&v�<(v�<4v�<v�<*v�<:v�<�u�<&v�<Dv�<v�<Dv�<&v�<�u�<:v�<*v�<v�<4v�<(v�<&v�<*v�<2v�<`   `   >v�<&v�<v�<�u�<Lv�<"v�<�u�< v�<2v�<�u�<�u�<;v�< v�<;v�<�u�<�u�<2v�< v�<�u�<"v�<Lv�<�u�<v�<&v�<`   `   �u�<v�<�u�<�u�<Pv�<v�<v�<�u�<�u�<8v�<	v�<6v�<v�<6v�<	v�<8v�<�u�<�u�<v�<v�<Pv�<�u�<�u�<v�<`   `   v�<>v�<(v�<#v�<Fv�<v�<Vv�<�u�<v�<Iv�<v�<,v�<v�<,v�<v�<Iv�<v�<�u�<Vv�<v�<Fv�<#v�<(v�<>v�<`   `   !v�<Ev�<v�<v�<9v�<v�<2v�<	v�<v�<*v�<v�<<v�<:v�<<v�<v�<*v�<v�<	v�<2v�<v�<9v�<v�<v�<Ev�<`   `   �u�<.v�<*v�<�u�<:v�<?v�<v�<v�<*v�<9v�<2v�< v�<=v�< v�<2v�<9v�<*v�<v�<v�<?v�<:v�<�u�<*v�<.v�<`   `   �u�<Iv�<Tv�<v�<v�< v�<,v�<?v�<.v�<+v�<*v�<�u�<v�<�u�<*v�<+v�<.v�<?v�<,v�< v�<v�<v�<Tv�<Iv�<`   `   �u�<v�<!v�<;v�<v�<�u�<v�<v�<v�<v�<0v�<>v�</v�<>v�<0v�<v�<v�<v�<v�<�u�<v�<;v�<!v�<v�<`   `   v�<�u�<�u�<@v�<7v�<v�<v�<v�<Jv�<Iv�<Bv�<Qv�<v�<Qv�<Bv�<Iv�<Jv�<v�<v�<v�<7v�<@v�<�u�<�u�<`   `   yv�<8v�<2v�<v�<v�<6v�<v�<v�<Cv�<Cv�<v�<)v�<v�<)v�<v�<Cv�<Cv�<v�<v�<6v�<v�<v�<2v�<8v�<`   `   Fv�<v�<_v�<v�<v�<av�<v�<v�<v�<v�<�u�<6v�<fv�<6v�<�u�<v�<v�<v�<v�<av�<v�<v�<_v�<v�<`   `   v�<�u�<5v�<v�<'v�<Qv�<.v�<av�< v�<v�<v�<v�<Ov�<v�<v�<v�< v�<av�<.v�<Qv�<'v�<v�<5v�<�u�<`   `   Lv�<&v�<�u�<�u�<v�<	v�<+v�<cv�<�u�<v�<#v�<�u�<Gv�<�u�<#v�<v�<�u�<cv�<+v�<	v�<v�<�u�<�u�<&v�<`   `   %v�<9v�<v�<
v�<+v�<v�<v�<-v�<�u�<>v�<@v�<v�<�v�<v�<@v�<>v�<�u�<-v�<v�<v�<+v�<
v�<v�<9v�<`   `   v�<.v�<4v�<+v�<'v�<_v�<5v�<v�<v�<9v�<v�<v�<uv�<v�<v�<9v�<v�<v�<5v�<_v�<'v�<+v�<4v�<.v�<`   `   Tv�<-v�<v�<v�<v�<jv�<Nv�<�u�<v�<�u�<v�<?v�<av�<?v�<v�<�u�<v�<�u�<Nv�<jv�<v�<v�<v�<-v�<`   `   �u�<v�<�u�<@v�<"v�<.v�<Bv�<v�<+v�<v�<^v�<uv�<5v�<uv�<^v�<v�<+v�<v�<Bv�<.v�<"v�<@v�<�u�<v�<`   `   �u�<v�<
v�<Gv�<5v�<v�<Vv�<v�<_v�<Fv�<v�<v�<�u�<v�<v�<Fv�<_v�<v�<Vv�<v�<5v�<Gv�<
v�<v�<`   `   0v�<]v�<,v�<"v�<v�<%v�<Wv�<v�<Gv�<0v�<�u�</v�<6v�</v�<�u�<0v�<Gv�<v�<Wv�<%v�<v�<"v�<,v�<]v�<`   `   v�<)v�<,v�<v�<v�<v�<.v�<5v�<v�<v�<v�<Rv�<Yv�<Rv�<v�<v�<v�<5v�<.v�<v�<v�<v�<,v�<)v�<`   `   �u�< v�<)v�<v�<8v�<�u�<v�<av�<v�<�u�<�u�<�u�<�u�<�u�<�u�<�u�<v�<av�<v�<�u�<8v�<v�<)v�< v�<`   `   Tv�<Dv�<;v�<v�<-v�<v�<v�<2v�<>v�<Mv�<
v�<%v�<+v�<%v�<
v�<Mv�<>v�<2v�<v�<v�<-v�<v�<;v�<Dv�<`   `   2v�< v�<<v�<"v�<v�<)v�<Mv�<v�<8v�<gv�<v�<Cv�<_v�<Cv�<v�<gv�<8v�<v�<Mv�<)v�<v�<"v�<<v�< v�<`   `   `v�<Fv�<Uv�<yv�<wv�<@v�<Sv�<iv�<7v�</v�<Mv�<Mv�< v�<Mv�<Mv�</v�<7v�<iv�<Sv�<@v�<wv�<yv�<Uv�<Fv�<`   `   Xv�<Lv�<Iv�<Sv�<ev�<Jv�<'v�<Pv�<:v�<Tv�<pv�<*v�<v�<*v�<pv�<Tv�<:v�<Pv�<'v�<Jv�<ev�<Sv�<Iv�<Lv�<`   `   4v�<Rv�<Sv�<@v�<Av�<hv�<Tv�<Xv�<Cv�<Tv�<wv�<Kv�<iv�<Kv�<wv�<Tv�<Cv�<Xv�<Tv�<hv�<Av�<@v�<Sv�<Rv�<`   `   v�<Xv�<kv�<Yv�<Hv�<�v�<�v�<\v�<Iv�<3v�<hv�<Rv�<[v�<Rv�<hv�<3v�<Iv�<\v�<�v�<�v�<Hv�<Yv�<kv�<Xv�<`   `   2v�<jv�<iv�<fv�<dv�<�v�<1v�<v�<Vv�<Mv�<Zv�<6v�<7v�<6v�<Zv�<Mv�<Vv�<v�<1v�<�v�<dv�<fv�<iv�<jv�<`   `   Nv�<Hv�<6v�<;v�<6v�<xv�<Av�<v�<Zv�<[v�<Iv�<?v�<xv�<?v�<Iv�<[v�<Zv�<v�<Av�<xv�<6v�<;v�<6v�<Hv�<`   `   Pv�<v�<&v�<Ev�<v�<Zv�<hv�<Wv�<Jv�<Nv�<Jv�<;v�<}v�<;v�<Jv�<Nv�<Jv�<Wv�<hv�<Zv�<v�<Ev�<&v�<v�<`   `   v�<Xv�<ev�<�v�<Ov�<Fv�<4v�<Jv�<Uv�<Mv�<Ev�<@v�<zv�<@v�<Ev�<Mv�<Uv�<Jv�<4v�<Fv�<Ov�<�v�<ev�<Xv�<`   `   Cv�<Dv�<6v�<Kv�<<v�<Nv�<Qv�<Uv�<ev�<Lv�<>v�<Xv�<�v�<Xv�<>v�<Lv�<ev�<Uv�<Qv�<Nv�<<v�<Kv�<6v�<Dv�<`   `   (v�<v�<�u�<6v�<(v�<Zv�<�v�<Nv�<;v�<Lv�<hv�<Sv�<rv�<Sv�<hv�<Lv�<;v�<Nv�<�v�<Zv�<(v�<6v�<�u�<v�<`   `   sv�<dv�<;v�<pv�<<v�<Kv�<Qv�<>v�<Jv�<Mv�<nv�<2v�<Ev�<2v�<nv�<Mv�<Jv�<>v�<Qv�<Kv�<<v�<pv�<;v�<dv�<`   `   v�<[v�<nv�<Vv�<v�<Gv�<v�<5v�<sv�<;v�<Dv�<%v�<Qv�<%v�<Dv�<;v�<sv�<5v�<v�<Gv�<v�<Vv�<nv�<[v�<`   `   �u�<Gv�<ov�<Pv�<2v�<nv�<;v�<v�<Wv�<<v�<\v�<Kv�<Yv�<Kv�<\v�<<v�<Wv�<v�<;v�<nv�<2v�<Pv�<ov�<Gv�<`   `   Bv�<fv�<=v�<`v�<_v�<Yv�<av�<;v�<rv�<`v�<dv�<hv�<[v�<hv�<dv�<`v�<rv�<;v�<av�<Yv�<_v�<`v�<=v�<fv�<`   `   ;v�<Yv�<2v�<Yv�<hv�<!v�<Av�<?v�<wv�<ev�<6v�<Kv�<:v�<Kv�<6v�<ev�<wv�<?v�<Av�<!v�<hv�<Yv�<2v�<Yv�<`   `   �u�<>v�<Wv�<Fv�<kv�<8v�<4v�< v�<3v�<Yv�<Lv�<@v�<�u�<@v�<Lv�<Yv�<3v�< v�<4v�<8v�<kv�<Fv�<Wv�<>v�<`   `   v�<v�<Vv�<Gv�<wv�<mv�<Cv�<8v�<;v�<Ov�<cv�<nv�<v�<nv�<cv�<Ov�<;v�<8v�<Cv�<mv�<wv�<Gv�<Vv�<v�<`   `   Ev�<#v�<cv�<Cv�<[v�<pv�<v�<&v�<bv�<Gv�<9v�<�v�<rv�<�v�<9v�<Gv�<bv�<&v�<v�<pv�<[v�<Cv�<cv�<#v�<`   `   iv�<Mv�<^v�<�u�<v�<fv�<v�<3v�<hv�<Tv�<5v�<iv�<pv�<iv�<5v�<Tv�<hv�<3v�<v�<fv�<v�<�u�<^v�<Mv�<`   `   Ev�<Av�<Uv�<$v�<Lv�<Zv�<-v�<bv�<8v�<1v�<Nv�<Bv�<<v�<Bv�<Nv�<1v�<8v�<bv�<-v�<Zv�<Lv�<$v�<Uv�<Av�<`   `   9v�<<v�<pv�<�v�<lv�<1v�<'v�<cv�<,v�<$v�<nv�<Nv�<7v�<Nv�<nv�<$v�<,v�<cv�<'v�<1v�<lv�<�v�<pv�<<v�<`   `   cv�<Rv�<Tv�<uv�<v�<%v�<`v�<kv�<wv�<Nv�<mv�<hv�<[v�<hv�<mv�<Nv�<wv�<kv�<`v�<%v�<v�<uv�<Tv�<Rv�<`   `   Xv�<Qv�<,v�<_v�<v�<0v�<dv�<1v�<jv�<2v�<v�<Cv�<_v�<Cv�<v�<2v�<jv�<1v�<dv�<0v�<v�<_v�<,v�<Qv�<`   `   Dv�<^v�<1v�<Qv�<@v�<Gv�<Kv�<v�<Pv�<Ev�<v�<.v�<Vv�<.v�<v�<Ev�<Pv�<v�<Kv�<Gv�<@v�<Qv�<1v�<^v�<`   `    v�<Mv�<Mv�</v�<7v�<iv�<Sv�<@v�<wv�<yv�<Uv�<Fv�<`v�<Fv�<Uv�<yv�<wv�<@v�<Sv�<iv�<7v�</v�<Mv�<Mv�<`   `   v�<*v�<pv�<Tv�<:v�<Pv�<'v�<Jv�<ev�<Sv�<Iv�<Lv�<Xv�<Lv�<Iv�<Sv�<ev�<Jv�<'v�<Pv�<:v�<Tv�<pv�<*v�<`   `   iv�<Kv�<wv�<Tv�<Cv�<Xv�<Tv�<hv�<Av�<@v�<Sv�<Rv�<4v�<Rv�<Sv�<@v�<Av�<hv�<Tv�<Xv�<Cv�<Tv�<wv�<Kv�<`   `   [v�<Rv�<hv�<3v�<Iv�<\v�<�v�<�v�<Hv�<Yv�<kv�<Xv�<v�<Xv�<kv�<Yv�<Hv�<�v�<�v�<\v�<Iv�<3v�<hv�<Rv�<`   `   7v�<6v�<Zv�<Mv�<Vv�<v�<1v�<�v�<dv�<fv�<iv�<jv�<2v�<jv�<iv�<fv�<dv�<�v�<1v�<v�<Vv�<Mv�<Zv�<6v�<`   `   xv�<?v�<Iv�<[v�<Zv�<v�<Av�<xv�<6v�<;v�<6v�<Hv�<Nv�<Hv�<6v�<;v�<6v�<xv�<Av�<v�<Zv�<[v�<Iv�<?v�<`   `   }v�<;v�<Jv�<Nv�<Jv�<Wv�<hv�<Zv�<v�<Ev�<&v�<v�<Pv�<v�<&v�<Ev�<v�<Zv�<hv�<Wv�<Jv�<Nv�<Jv�<;v�<`   `   zv�<@v�<Ev�<Mv�<Uv�<Jv�<4v�<Fv�<Ov�<�v�<ev�<Xv�<v�<Xv�<ev�<�v�<Ov�<Fv�<4v�<Jv�<Uv�<Mv�<Ev�<@v�<`   `   �v�<Xv�<>v�<Lv�<ev�<Uv�<Qv�<Nv�<<v�<Kv�<6v�<Dv�<Cv�<Dv�<6v�<Kv�<<v�<Nv�<Qv�<Uv�<ev�<Lv�<>v�<Xv�<`   `   rv�<Sv�<hv�<Lv�<;v�<Nv�<�v�<Zv�<(v�<6v�<�u�<v�<(v�<v�<�u�<6v�<(v�<Zv�<�v�<Nv�<;v�<Lv�<hv�<Sv�<`   `   Ev�<2v�<nv�<Mv�<Jv�<>v�<Qv�<Kv�<<v�<pv�<;v�<dv�<sv�<dv�<;v�<pv�<<v�<Kv�<Qv�<>v�<Jv�<Mv�<nv�<2v�<`   `   Qv�<%v�<Dv�<;v�<sv�<5v�<v�<Gv�<v�<Vv�<nv�<[v�<v�<[v�<nv�<Vv�<v�<Gv�<v�<5v�<sv�<;v�<Dv�<%v�<`   `   Yv�<Kv�<\v�<<v�<Wv�<v�<;v�<nv�<2v�<Pv�<ov�<Gv�<�u�<Gv�<ov�<Pv�<2v�<nv�<;v�<v�<Wv�<<v�<\v�<Kv�<`   `   [v�<hv�<dv�<`v�<rv�<;v�<av�<Yv�<_v�<`v�<=v�<fv�<Bv�<fv�<=v�<`v�<_v�<Yv�<av�<;v�<rv�<`v�<dv�<hv�<`   `   :v�<Kv�<6v�<ev�<wv�<?v�<Av�<!v�<hv�<Yv�<2v�<Yv�<;v�<Yv�<2v�<Yv�<hv�<!v�<Av�<?v�<wv�<ev�<6v�<Kv�<`   `   �u�<@v�<Lv�<Yv�<3v�< v�<4v�<8v�<kv�<Fv�<Wv�<>v�<�u�<>v�<Wv�<Fv�<kv�<8v�<4v�< v�<3v�<Yv�<Lv�<@v�<`   `   v�<nv�<cv�<Ov�<;v�<8v�<Cv�<mv�<wv�<Gv�<Vv�<v�<v�<v�<Vv�<Gv�<wv�<mv�<Cv�<8v�<;v�<Ov�<cv�<nv�<`   `   rv�<�v�<9v�<Gv�<bv�<&v�<v�<pv�<[v�<Cv�<cv�<#v�<Ev�<#v�<cv�<Cv�<[v�<pv�<v�<&v�<bv�<Gv�<9v�<�v�<`   `   pv�<iv�<5v�<Tv�<hv�<3v�<v�<fv�<v�<�u�<^v�<Mv�<iv�<Mv�<^v�<�u�<v�<fv�<v�<3v�<hv�<Tv�<5v�<iv�<`   `   <v�<Bv�<Nv�<1v�<8v�<bv�<-v�<Zv�<Lv�<$v�<Uv�<Av�<Ev�<Av�<Uv�<$v�<Lv�<Zv�<-v�<bv�<8v�<1v�<Nv�<Bv�<`   `   7v�<Nv�<nv�<$v�<,v�<cv�<'v�<1v�<lv�<�v�<pv�<<v�<9v�<<v�<pv�<�v�<lv�<1v�<'v�<cv�<,v�<$v�<nv�<Nv�<`   `   [v�<hv�<mv�<Nv�<wv�<kv�<`v�<%v�<v�<uv�<Tv�<Rv�<cv�<Rv�<Tv�<uv�<v�<%v�<`v�<kv�<wv�<Nv�<mv�<hv�<`   `   _v�<Cv�<v�<2v�<jv�<1v�<dv�<0v�<v�<_v�<,v�<Qv�<Xv�<Qv�<,v�<_v�<v�<0v�<dv�<1v�<jv�<2v�<v�<Cv�<`   `   Vv�<.v�<v�<Ev�<Pv�<v�<Kv�<Gv�<@v�<Qv�<1v�<^v�<Dv�<^v�<1v�<Qv�<@v�<Gv�<Kv�<v�<Pv�<Ev�<v�<.v�<`   `   �v�<�v�<nv�<Hv�<Vv�<�v�<}v�<rv�<�v�<rv�<�v�<�v�<�v�<�v�<�v�<rv�<�v�<rv�<}v�<�v�<Vv�<Hv�<nv�<�v�<`   `   �v�<Lv�<jv�<�v�<=v�<|v�<�v�<yv�<�v�<�v�<\v�<qv�<�v�<qv�<\v�<�v�<�v�<yv�<�v�<|v�<=v�<�v�<jv�<Lv�<`   `   �v�<tv�<�v�<�v�<pv�<fv�<�v�<hv�<`v�<�v�<dv�<Qv�<�v�<Qv�<dv�<�v�<`v�<hv�<�v�<fv�<pv�<�v�<�v�<tv�<`   `   �v�<nv�<Jv�<ev�<{v�<dv�<fv�<�v�<ev�<�v�<�v�<vv�<�v�<vv�<�v�<�v�<ev�<�v�<fv�<dv�<{v�<ev�<Jv�<nv�<`   `   �v�<pv�<Fv�<Fv�<xv�<Mv�<@v�<�v�<|v�<gv�<�v�<iv�<�v�<iv�<�v�<gv�<|v�<�v�<@v�<Mv�<xv�<Fv�<Fv�<pv�<`   `   ov�<�v�<�v�<�v�<�v�<xv�<wv�<�v�<rv�<kv�<�v�<^v�<�v�<^v�<�v�<kv�<rv�<�v�<wv�<xv�<�v�<�v�<�v�<�v�<`   `   dv�<�v�<�v�<�v�<�v�<v�<�v�<{v�<Ov�<�v�<�v�<av�<�v�<av�<�v�<�v�<Ov�<{v�<�v�<v�<�v�<�v�<�v�<�v�<`   `   wv�<�v�<cv�<Sv�<�v�<{v�<av�<wv�<rv�<�v�<�v�<Jv�<�v�<Jv�<�v�<�v�<rv�<wv�<av�<{v�<�v�<Sv�<cv�<�v�<`   `   `v�<�v�<�v�<}v�<�v�<�v�<sv�<�v�<�v�<Zv�<|v�<pv�<uv�<pv�<|v�<Zv�<�v�<�v�<sv�<�v�<�v�<}v�<�v�<�v�<`   `   yv�<�v�<�v�<�v�<ov�<iv�<Yv�<{v�<rv�<Tv�<�v�<�v�<_v�<�v�<�v�<Tv�<rv�<{v�<Yv�<iv�<ov�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<zv�<qv�<�v�<�v�<{v�<jv�<Nv�<jv�<{v�<�v�<�v�<qv�<zv�<�v�<�v�<�v�<�v�<�v�<`   `   jv�<qv�<Ov�<wv�<�v�<�v�<�v�<�v�<�v�<{v�<]v�<�v�<�v�<�v�<]v�<{v�<�v�<�v�<�v�<�v�<�v�<wv�<Ov�<qv�<`   `   �v�<�v�<^v�<�v�<�v�<Dv�<�v�<vv�<jv�<nv�<�v�<�v�<�v�<�v�<�v�<nv�<jv�<vv�<�v�<Dv�<�v�<�v�<^v�<�v�<`   `   �v�<�v�<Qv�<�v�<�v�<v�<�v�<�v�<pv�<�v�<�v�<Uv�<(v�<Uv�<�v�<�v�<pv�<�v�<�v�<v�<�v�<�v�<Qv�<�v�<`   `   v�<�v�<Yv�<[v�<�v�<}v�<�v�<�v�<`v�<kv�<iv�<�v�<�v�<�v�<iv�<kv�<`v�<�v�<�v�<}v�<�v�<[v�<Yv�<�v�<`   `   zv�<�v�<�v�<Hv�<pv�<�v�<�v�<nv�<wv�<wv�<]v�<�v�<�v�<�v�<]v�<wv�<wv�<nv�<�v�<�v�<pv�<Hv�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<Tv�<hv�<�v�<�v�<�v�<�v�<sv�<iv�<Mv�<iv�<sv�<�v�<�v�<�v�<�v�<hv�<Tv�<�v�<�v�<�v�<`   `   �v�< v�<Mv�<�v�<ov�<pv�<�v�<�v�<kv�<]v�<�v�<jv�<Bv�<jv�<�v�<]v�<kv�<�v�<�v�<pv�<ov�<�v�<Mv�< v�<`   `   �v�<vv�<�v�<�v�<lv�<�v�<�v�<�v�<Kv�<vv�<�v�<{v�<�v�<{v�<�v�<vv�<Kv�<�v�<�v�<�v�<lv�<�v�<�v�<vv�<`   `   �v�<rv�<�v�<|v�<sv�<�v�<}v�<�v�<�v�<�v�<�v�<Ev�<�v�<Ev�<�v�<�v�<�v�<�v�<}v�<�v�<sv�<|v�<�v�<rv�<`   `   `v�<Tv�<Nv�<Wv�<v�<�v�<pv�<�v�<�v�<�v�<Vv�<Tv�<�v�<Tv�<Vv�<�v�<�v�<�v�<pv�<�v�<v�<Wv�<Nv�<Tv�<`   `   �v�<�v�<xv�<fv�<�v�<�v�<�v�<dv�<[v�<�v�<pv�<vv�<�v�<vv�<pv�<�v�<[v�<dv�<�v�<�v�<�v�<fv�<xv�<�v�<`   `   8v�<�v�<�v�<qv�<�v�<�v�<�v�<�v�<tv�<�v�<�v�<kv�<7v�<kv�<�v�<�v�<tv�<�v�<�v�<�v�<�v�<qv�<�v�<�v�<`   `   v�<{v�<�v�<hv�<�v�<jv�<]v�<�v�<�v�<|v�<�v�<�v�<mv�<�v�<�v�<|v�<�v�<�v�<]v�<jv�<�v�<hv�<�v�<{v�<`   `   �v�<�v�<�v�<rv�<�v�<rv�<}v�<�v�<Vv�<Hv�<nv�<�v�<�v�<�v�<nv�<Hv�<Vv�<�v�<}v�<rv�<�v�<rv�<�v�<�v�<`   `   �v�<qv�<\v�<�v�<�v�<yv�<�v�<|v�<=v�<�v�<jv�<Lv�<�v�<Lv�<jv�<�v�<=v�<|v�<�v�<yv�<�v�<�v�<\v�<qv�<`   `   �v�<Qv�<dv�<�v�<`v�<hv�<�v�<fv�<pv�<�v�<�v�<tv�<�v�<tv�<�v�<�v�<pv�<fv�<�v�<hv�<`v�<�v�<dv�<Qv�<`   `   �v�<vv�<�v�<�v�<ev�<�v�<fv�<dv�<{v�<ev�<Jv�<nv�<�v�<nv�<Jv�<ev�<{v�<dv�<fv�<�v�<ev�<�v�<�v�<vv�<`   `   �v�<iv�<�v�<gv�<|v�<�v�<@v�<Mv�<xv�<Fv�<Fv�<pv�<�v�<pv�<Fv�<Fv�<xv�<Mv�<@v�<�v�<|v�<gv�<�v�<iv�<`   `   �v�<^v�<�v�<kv�<rv�<�v�<wv�<xv�<�v�<�v�<�v�<�v�<ov�<�v�<�v�<�v�<�v�<xv�<wv�<�v�<rv�<kv�<�v�<^v�<`   `   �v�<av�<�v�<�v�<Ov�<{v�<�v�<v�<�v�<�v�<�v�<�v�<dv�<�v�<�v�<�v�<�v�<v�<�v�<{v�<Ov�<�v�<�v�<av�<`   `   �v�<Jv�<�v�<�v�<rv�<wv�<av�<{v�<�v�<Sv�<cv�<�v�<wv�<�v�<cv�<Sv�<�v�<{v�<av�<wv�<rv�<�v�<�v�<Jv�<`   `   uv�<pv�<|v�<Zv�<�v�<�v�<sv�<�v�<�v�<}v�<�v�<�v�<`v�<�v�<�v�<}v�<�v�<�v�<sv�<�v�<�v�<Zv�<|v�<pv�<`   `   _v�<�v�<�v�<Tv�<rv�<{v�<Yv�<iv�<ov�<�v�<�v�<�v�<yv�<�v�<�v�<�v�<ov�<iv�<Yv�<{v�<rv�<Tv�<�v�<�v�<`   `   Nv�<jv�<{v�<�v�<�v�<qv�<zv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<zv�<qv�<�v�<�v�<{v�<jv�<`   `   �v�<�v�<]v�<{v�<�v�<�v�<�v�<�v�<�v�<wv�<Ov�<qv�<jv�<qv�<Ov�<wv�<�v�<�v�<�v�<�v�<�v�<{v�<]v�<�v�<`   `   �v�<�v�<�v�<nv�<jv�<vv�<�v�<Dv�<�v�<�v�<^v�<�v�<�v�<�v�<^v�<�v�<�v�<Dv�<�v�<vv�<jv�<nv�<�v�<�v�<`   `   (v�<Uv�<�v�<�v�<pv�<�v�<�v�<v�<�v�<�v�<Qv�<�v�<�v�<�v�<Qv�<�v�<�v�<v�<�v�<�v�<pv�<�v�<�v�<Uv�<`   `   �v�<�v�<iv�<kv�<`v�<�v�<�v�<}v�<�v�<[v�<Yv�<�v�<v�<�v�<Yv�<[v�<�v�<}v�<�v�<�v�<`v�<kv�<iv�<�v�<`   `   �v�<�v�<]v�<wv�<wv�<nv�<�v�<�v�<pv�<Hv�<�v�<�v�<zv�<�v�<�v�<Hv�<pv�<�v�<�v�<nv�<wv�<wv�<]v�<�v�<`   `   Mv�<iv�<sv�<�v�<�v�<�v�<�v�<hv�<Tv�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<Tv�<hv�<�v�<�v�<�v�<�v�<sv�<iv�<`   `   Bv�<jv�<�v�<]v�<kv�<�v�<�v�<pv�<ov�<�v�<Mv�< v�<�v�< v�<Mv�<�v�<ov�<pv�<�v�<�v�<kv�<]v�<�v�<jv�<`   `   �v�<{v�<�v�<vv�<Kv�<�v�<�v�<�v�<lv�<�v�<�v�<vv�<�v�<vv�<�v�<�v�<lv�<�v�<�v�<�v�<Kv�<vv�<�v�<{v�<`   `   �v�<Ev�<�v�<�v�<�v�<�v�<}v�<�v�<sv�<|v�<�v�<rv�<�v�<rv�<�v�<|v�<sv�<�v�<}v�<�v�<�v�<�v�<�v�<Ev�<`   `   �v�<Tv�<Vv�<�v�<�v�<�v�<pv�<�v�<v�<Wv�<Nv�<Tv�<`v�<Tv�<Nv�<Wv�<v�<�v�<pv�<�v�<�v�<�v�<Vv�<Tv�<`   `   �v�<vv�<pv�<�v�<[v�<dv�<�v�<�v�<�v�<fv�<xv�<�v�<�v�<�v�<xv�<fv�<�v�<�v�<�v�<dv�<[v�<�v�<pv�<vv�<`   `   7v�<kv�<�v�<�v�<tv�<�v�<�v�<�v�<�v�<qv�<�v�<�v�<8v�<�v�<�v�<qv�<�v�<�v�<�v�<�v�<tv�<�v�<�v�<kv�<`   `   mv�<�v�<�v�<|v�<�v�<�v�<]v�<jv�<�v�<hv�<�v�<{v�<v�<{v�<�v�<hv�<�v�<jv�<]v�<�v�<�v�<|v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   %w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   `   �v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<%w�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<�v�<`   