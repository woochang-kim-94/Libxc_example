H   �0�ŀ�@                }�ŀ�@ �,Gܞ@                        rdB �G@H            �         `   c��<���<���<E��<R��<���<e��<a��<���<���<���<u��<l��<u��<���<���<���<a��<>��<���<t��<E��<���<���<`   `   ���<H��<J��<{��<-��<G��<���<̆�<���<R��<U��<|��<q��<U��<f��<���<���<���<^��<��<j��<V��<O��<~��<`   `   ���<J��<h��<r��<}��<���<��<���<���<U��<��<%��<$��<U��<���<���< ��<���<v��<r��<n��<J��<���<��<`   `   E��<{��<r��<��<8��<m��<b��<]��<k��<���<���<���<���<a��<q��<r��<T��<'��<
��<~��<j��<B��<~��<w��<`   `   R��<-��<}��<8��<:��<���<���<E��<}��<S��<J��<S��<���<E��<~��<���<c��<8��<Y��<-��<f��<!��<D��<!��<`   `   ���<G��<���<m��<���<_��<.��<���<y��<M��<M��<p��<���<>��<s��<���<T��<���<^��<���<���<]��<e��<���<`   `   e��<���<��<b��<���<.��<Y��<Ć�<���<���<���<Ć�<U��<.��<���<b��<$��<���<Q��<���<w��<���<_��<���<`   `   a��<̆�<���<]��<E��<���<Ć�<T��<R��<I��<U��<ӆ�<���<4��<q��<���<���<^��<��<��<J��<\��<&��<���<`   `   ���<���<���<k��<}��<y��<���<R��<_��<R��<z��<y��<���<k��<r��<���<���<`��<W��< ��<!��< ��<g��<`��<`   `   ���<R��<U��<���<S��<M��<���<I��<R��<ʆ�<M��<C��<���<a��<f��<���<��<���<b��<���<���<K��<���<���<`   `   ���<U��<��<���<J��<M��<���<U��<z��<M��<Z��<���<��<U��<���< ��<7��<���<T��<=��<|��<���<��< ��<`   `   u��<|��<%��<���<S��<p��<Ć�<ӆ�<y��<C��<���<1��<q��<r��<9��<C��<5��<M��<��<���<;��<N��<J��<%��<`   `   l��<q��<$��<���<���<���<U��<���<���<���<��<q��<z��<(��<���<���<	��<q��<���<q��<��<���<Ɔ�<(��<`   `   u��<U��<U��<a��<E��<>��<.��<4��<k��<a��<U��<r��<(��<��<1��<���<w��< ��<��<���<��<��<&��<3��<`   `   ���<f��<���<q��<~��<s��<���<q��<r��<f��<���<9��<���<1��<-��<h��<g��<��<8��<h��<R��<1��<���<9��<`   `   ���<���<���<r��<���<���<b��<���<���<���< ��<C��<���<���<h��<N��<w��<���<e��<T��<��<���<J��< ��<`   `   ���<���< ��<T��<c��<T��<$��<���<���<��<7��<5��<	��<w��<g��<w��<��<w��<d��<w��<��<5��<0��<��<`   `   a��<���<���<'��<8��<���<���<^��<`��<���<���<M��<q��< ��<��<���<w��<��<��<|��<;��<���<���<W��<`   `   >��<^��<v��<
��<Y��<^��<Q��<��<W��<b��<T��<��<���<��<8��<e��<d��<��<���<��<e��<b��<Y��<��<`   `   ���<��<r��<~��<-��<���<���<��< ��<���<=��<���<q��<���<h��<T��<w��<|��<��<=��<���<��<&��<���<`   `   t��<j��<n��<j��<f��<���<w��<J��<!��<���<|��<;��<��<��<R��<��<��<;��<e��<���<<��<J��<`��<���<`   `   E��<V��<J��<B��<!��<]��<���<\��< ��<K��<���<N��<���<��<1��<���<5��<���<b��<��<J��<���<e��<��<`   `   ���<O��<���<~��<D��<e��<_��<&��<g��<���<��<J��<Ɔ�<&��<���<J��<0��<���<Y��<&��<`��<e��<M��<~��<`   `   ���<~��<��<w��<!��<���<���<���<`��<���< ��<%��<(��<3��<9��< ��<��<W��<��<���<���<��<~��<��<`   `   ���<L��<a��<���<u��<k��<���<q��<��<V��<���<h��<h��<h��<���<V��<=��<q��<j��<k��<���<���<N��<L��<`   `   L��<p��<���<���<c��<5��<b��<t��<)��<@��<u��<���<���<u��<S��< ��<]��<r��<K��<R��<���<���<v��<I��<`   `   a��<���<=��<���<���<���<��<p��<���<���<c��<���<m��<���<w��<p��<��<���<���<���<B��<���<]��<��<`   `   ���<���<���<i��<���<���<x��<M��<T��<���<|��<|��<u��<K��<`��<���<���<|��<���<���<���<���<_��<X��<`   `   u��<c��<���<���<o��<M��<���<f��<R��<O��<���<O��<f��<f��<o��<M��<���<���<���<c��<���<v��<�<v��<`   `   k��<5��<���<���<M��<>��<���<���<J��<z��<{��<A��<v��<���<Q��<=��<���<���<K��<g��<[��<e��<l��<k��<`   `   ���<b��<��<x��<���<���<,��<>��<R��<j��<[��<>��<'��<���<���<x��<!��<b��<|��<v��<;��<r��<#��<v��<`   `   q��<t��<p��<M��<f��<���<>��<Q��<m��<d��<Q��<M��<v��<V��<`��<{��<]��<n��<���<���<���<���<���<���<`   `   ��<)��<���<T��<R��<J��<R��<m��<ņ�<m��<C��<J��<m��<T��<b��<)��<7��<m��<Ć�<���<i��<���<Ԇ�<m��<`   `   V��<@��<���<���<O��<z��<j��<d��<m��<z��<{��<?��<u��<���<S��<S��<~��<S��<@��<���<���<)��<Z��<���<`   `   ���<u��<c��<|��<���<{��<[��<Q��<C��<{��<���<|��<a��<u��<���<���<���<���<p��<���<���<���<r��<���<`   `   h��<���<���<|��<O��<A��<>��<M��<J��<?��<|��<���<���<e��<g��<v��<���<���<~��<h��<���<���<}��<T��<`   `   h��<���<m��<u��<f��<v��<'��<v��<m��<u��<a��<���<v��<���<���<o��<>��<���<ņ�<���<7��<o��<���<���<`   `   h��<u��<���<K��<f��<���<���<V��<T��<���<u��<e��<���<���<c��<���<���<c��<z��<���<���<O��<���<���<`   `   ���<S��<w��<`��<o��<Q��<���<`��<b��<S��<���<g��<���<c��<���<c��<���<���<w��<c��<���<c��<���<g��<`   `   V��< ��<p��<���<M��<=��<x��<{��<)��<S��<���<v��<o��<���<c��<7��<���<���<N��<P��<���<y��<}��<���<`   `   =��<]��<��<���<���<���<!��<]��<7��<~��<���<���<>��<���<���<���<��<���<���<���<D��<���<���<~��<`   `   q��<r��<���<|��<���<���<b��<n��<m��<S��<���<���<���<c��<���<���<���<���<z��<���<���<���<Z��<c��<`   `   j��<K��<���<���<���<K��<|��<���<Ć�<@��<p��<~��<ņ�<z��<w��<N��<���<z��<���<~��<���<@��<ǆ�<���<`   `   k��<R��<���<���<c��<g��<v��<���<���<���<���<h��<���<���<c��<P��<���<���<~��<���<���<���<���<���<`   `   ���<���<B��<���<���<[��<;��<���<i��<���<���<���<7��<���<���<���<D��<���<���<���<���<���<$��<[��<`   `   ���<���<���<���<v��<e��<r��<���<���<)��<���<���<o��<O��<c��<y��<���<���<@��<���<���<���<l��<f��<`   `   N��<v��<]��<_��<�<l��<#��<���<Ԇ�<Z��<r��<}��<���<���<���<}��<���<Z��<ǆ�<���<$��<l��<ˆ�<_��<`   `   L��<I��<��<X��<v��<k��<v��<���<m��<���<���<T��<���<���<g��<���<~��<c��<���<���<[��<f��<_��<$��<`   `   چ�<���<���<���<x��<���<���<���<���<���<���<d��<O��<d��<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<���<h��<���<ن�<���<|��<���<���<}��<���<���<���<Ć�<���<|��<���<���<���<���<���<`   `   ���<���<��<���<���<i��<l��<���<ņ�<���<{��<���<���<���<���<���<r��<i��<���<���<��<���<���<���<`   `   ���<���<���<Y��<W��<φ�<���<X��<���<���<\��<\��<w��<��<i��<ˆ�<���<H��<l��<���<���<���<���<~��<`   `   x��<���<���<W��<���<q��<���<���<���<���<���<���<���<���<x��<q��<���<W��<���<���<���<|��<���<|��<`   `   ���<h��<i��<φ�<q��<R��<Ć�<���<���<���<���<���<���<ӆ�<b��<b��<���<t��<|��<���<���<���<���<���<`   `   ���<���<l��<���<���<Ć�<L��<���<���<J��<���<���<G��<Ć�<���<���<u��<���<���<���<m��<���<Y��<���<`   `   ���<ن�<���<X��<���<���<���<���<���<w��<���<���<���<��<i��<ņ�<Ć�<���<\��<f��<���<���<l��<H��<`   `   ���<���<ņ�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<t��<���<���<6��<���<���<t��<`   `   ���<|��<���<���<���<���<J��<w��<���<X��<���<w��<w��<Æ�<���<���<���<Z��<f��<���<y��<R��<`��<���<`   `   ���<���<{��<\��<���<���<���<���<���<���<���<\��<y��<���<���<���<���<e��<x��<���<���<e��<k��<���<`   `   d��<���<���<\��<���<���<���<���<���<w��<\��<���<}��<`��<p��<e��<���<���<`��<M��<���<Æ�<j��<_��<`   `   O��<}��<���<w��<���<���<G��<���<���<w��<y��<}��<[��<���<]��<^��<Q��<c��<n��<c��<K��<^��<h��<���<`   `   d��<���<���<��<���<ӆ�<Ć�<��<���<Æ�<���<`��<���<���<z��<���<���<P��<d��<���<���<i��<���<���<`   `   ���<���<���<i��<x��<b��<���<i��<���<���<���<p��<]��<z��<���<i��<���<m��<y��<i��<چ�<z��<N��<p��<`   `   ���<���<���<ˆ�<q��<b��<���<ņ�<���<���<���<e��<^��<���<i��<O��<���<���<c��<X��<���<g��<j��<���<`   `   ���<Ć�<r��<���<���<���<u��<Ć�<���<���<���<���<Q��<���<���<���<%��<���<���<���<V��<���<��<���<`   `   ���<���<i��<H��<W��<t��<���<���<t��<Z��<e��<���<c��<P��<m��<���<���<\��<d��<l��<���<f��<`��<k��<`   `   ���<|��<���<l��<���<|��<���<\��<���<f��<x��<`��<n��<d��<y��<c��<���<d��<R��<`��<���<f��<���<\��<`   `   ���<���<���<���<���<���<���<f��<���<���<���<M��<c��<���<i��<X��<���<l��<`��<���<y��<y��<l��<���<`   `   ���<���<��<���<���<���<m��<���<6��<y��<���<���<K��<���<چ�<���<V��<���<���<y��<M��<���<Y��<���<`   `   ���<���<���<���<|��<���<���<���<���<R��<e��<Æ�<^��<i��<z��<g��<���<f��<f��<y��<���<���<���<l��<`   `   ���<���<���<���<���<���<Y��<l��<���<`��<k��<j��<h��<���<N��<j��<��<`��<���<l��<Y��<���<Ć�<���<`   `   ���<���<���<~��<|��<���<���<H��<t��<���<���<_��<���<���<p��<���<���<k��<\��<���<���<l��<���<���<`   `   f��<���<���<���<���<���<ӆ�<���<���<���<ֆ�<��<���<��<ǆ�<���<Ɔ�<���<���<���<���<���<���<���<`   `   ���<e��<ˆ�<��<���<���<̆�<���<���<���<���<ц�<ʆ�<���<���<���<���<ن�<���<���<��<ֆ�<i��<���<`   `   ���<ˆ�<Ć�<׆�<���<҆�<b��<���<���<���<���<܆�<���<���<���<���<f��<҆�<���<׆�<ņ�<ˆ�<���<��<`   `   ���<��<׆�<���<���<׆�<���<���<���<ӆ�<Ά�<φ�<͆�<���<���<Ć�<ǆ�<���<���<��<��<���<�<���<`   `   ���<���<���<���<���<Ɔ�<���<���<ӆ�<���<���<���<��<���<Ɔ�<Ɔ�<φ�<���<߆�<���<���<���<���<���<`   `   ���<���<҆�<׆�<Ɔ�<���<���<���<���<���<���<���<���<���<Ɔ�<���<ǆ�<݆�<���<���<��<���<���<��<`   `   ӆ�<̆�<b��<���<���<���<���<Ȇ�<���<��<���<Ȇ�<���<���<���<���<h��<̆�<ǆ�<���<��<̆�<���<���<`   `   ���<���<���<���<���<���<Ȇ�<���<���<���<���<Ն�<���<���<���<���<���<���<~��<���<І�<ۆ�<���<n��<`   `   ���<���<���<���<ӆ�<���<���<���<ʆ�<���<���<���<��<���<���<���<���<���<��<���<���<���<��<���<`   `   ���<���<���<ӆ�<���<���<��<���<���<���<���<���<͆�<���<���<���<̆�<��<��<��<߆�<��<���<݆�<`   `   ֆ�<���<���<Ά�<���<���<���<���<���<���<���<Ά�<���<���<͆�<���<���<���<���<���<ۆ�<���<x��<���<`   `   ��<ц�<܆�<φ�<���<���<Ȇ�<Ն�<���<���<Ά�<��<ʆ�<��<Ն�<͆�<ކ�<���<���<���<���<��<ц�<Ȇ�<`   `   ���<ʆ�<���<͆�<��<���<���<���<��<͆�<���<ʆ�<���<�<ۆ�<	��<���<ކ�</��<ކ�<���<	��<��<�<`   `   ��<���<���<���<���<���<���<���<���<���<���<��<�<���<Ɔ�<ʆ�<��<̆�<ۆ�<���<���<���<���<Ɇ�<`   `   ǆ�<���<���<���<Ɔ�<Ɔ�<���<���<���<���<͆�<Ն�<ۆ�<Ɔ�<���<���<��<d��<҆�<���<���<Ɔ�<ц�<Ն�<`   `   ���<���<���<Ć�<Ɔ�<���<���<���<���<���<���<͆�<	��<ʆ�<���<��<؆�<��<��<���<���<��<ц�<���<`   `   Ɔ�<���<f��<ǆ�<φ�<ǆ�<h��<���<���<̆�<���<ކ�<���<��<��<؆�<ˆ�<؆�<���<��<���<ކ�<���<̆�<`   `   ���<ن�<҆�<���<���<݆�<̆�<���<���<��<���<���<ކ�<̆�<d��<��<؆�<W��<ۆ�<��<���<���<���<���<`   `   ���<���<���<���<߆�<���<ǆ�<~��<��<��<���<���</��<ۆ�<҆�<��<���<ۆ�<��<���<ˆ�<��<��<~��<`   `   ���<���<׆�<��<���<���<���<���<���<��<���<���<ކ�<���<���<���<��<��<���<���<߆�<���<���<��<`   `   ���<��<ņ�<��<���<��<��<І�<���<߆�<ۆ�<���<���<���<���<���<���<���<ˆ�<߆�<Ɇ�<І�<ކ�<��<`   `   ���<ֆ�<ˆ�<���<���<���<̆�<ۆ�<���<��<���<��<	��<���<Ɔ�<��<ކ�<���<��<���<І�<ن�<���<���<`   `   ���<i��<���<�<���<���<���<���<��<���<x��<ц�<��<���<ц�<ц�<���<���<��<���<ކ�<���<���<�<`   `   ���<���<��<���<���<��<���<n��<���<݆�<���<Ȇ�<�<Ɇ�<Ն�<���<̆�<���<~��<��<��<���<�<)��<`   `   O��<(��<ۆ�<���<��<���<��<��<׆�<��<��<��<ӆ�<��<���<��<��<��<���<���<(��<���<ц�<(��<`   `   (��<+��<��<��<��<Ն�<��<��<	��<���<��<��<���<��<���<��<��<'��<߆�<��<	��<��<-��<#��<`   `   ۆ�<��<���<ц�<��<	��<��< ��<#��<���<ن�<��<ۆ�<���<"��< ��<��<	��<	��<ц�<���<��<ކ�<ֆ�<`   `   ���<��<ц�<ӆ�<��<��<	��<��<���<���<��<��<���<��<��<��<���<���<݆�<چ�<	��<���<��<��<`   `   ��<��<��<��<���<Ć�<)��<��<���<���<��<���<��<��<��<Ć�<��<��<��<��< ��<0��<W��<0��<`   `   ���<Ն�<	��<��<Ć�<��<��<��<���<���<���<��<	��<��<���<���<���<��<߆�<���<׆�<��<��<ކ�<`   `   ��<��<��<	��<)��<��<*��<1��<��<y��<���<1��<#��<��<,��<	��<��<��<��<���<���<͆�<���<���<`   `   ��<��< ��<��<��<��<1��<���<��<���<���<<��<	��<��<��<)��<��<���<;��<���<��<��<��<0��<`   `   ׆�<	��<#��<���<���<���<��<��<(��<��<��<���<��<���<��<	��<��<��<��<̆�<��<̆�<
��<��<`   `   ��<���<���<���<���<���<y��<���<��<���<���<��<���<��<���< ��<��<҆�<���<��<ކ�<���<ӆ�<��<`   `   ��<��<ن�<��<��<���<���<���<��<���<��<��<Ԇ�<��<��<��<���<��<��<ʆ�<���<��<��<��<`   `   ��<��<��<��<���<��<1��<<��<���<��<��<��<���<��<چ�<��<���<��<��<��<��<��<���<ц�<`   `   ӆ�<���<ۆ�<���<��<	��<#��<	��<��<���<Ԇ�<���<ۆ�<��<��<ن�<���<׆�<��<׆�<���<ن�<��<��<`   `   ��<��<���<��<��<��<��<��<���<��<��<��<��<���<���<���<���<Æ�<Ά�<���<��<��<���<��<`   `   ���<���<"��<��<��<���<,��<��<��<���<��<چ�<��<���<��<��<��<��<���<��<��<���<��<چ�<`   `   ��<��< ��<��<Ć�<���<	��<)��<	��< ��<��<��<ن�<���<��<���<��<��<�<��<��<݆�<���<��<`   `   ��<��<��<���<��<���<��<��<��<��<���<���<���<���<��<��<Ć�<��<��<���<���<���<��<��<`   `   ��<'��<	��<���<��<��<��<���<��<҆�<��<��<׆�<Æ�<��<��<��<��<Ά�<چ�<��<��<ӆ�<��<`   `   ���<߆�<	��<݆�<��<߆�<��<;��<��<���<��<��<��<Ά�<���<�<��<Ά�<׆�<��<��<���<��<;��<`   `   ���<��<ц�<چ�<��<���<���<���<̆�<��<ʆ�<��<׆�<���<��<��<���<چ�<��<̆�<ކ�<Ć�<��<��<`   `   (��<	��<���<	��< ��<׆�<���<��<��<ކ�<���<��<���<��<��<��<���<��<��<ކ�<&��<��<���<׆�<`   `   ���<��<��<���<0��<��<͆�<��<̆�<���<��<��<ن�<��<���<݆�<���<��<���<Ć�<��<؆�<��<$��<`   `   ц�<-��<ކ�<��<W��<��<���<��<
��<ӆ�<��<���<��<���<��<���<��<ӆ�<��<��<���<��<`��<��<`   `   (��<#��<ֆ�<��<0��<ކ�<���<0��<��<��<��<ц�<��<��<چ�<��<��<��<;��<��<׆�<$��<��<߆�<`   `   ��<$��<Y��<0��<Z��<���<C��<,��<M��<G��<5��<2��<j��<2��<.��<G��<X��<,��<6��<���<f��<0��<S��<$��<`   `   $��<`��<N��<4��<~��<U��<E��<o��<8��<2��<^��<g��<g��<a��<6��<2��<j��<M��<Z��<u��<2��<U��<`��< ��<`   `   Y��<N��<,��<���<K��<��<>��<8��<3��<j��<S��<Q��<Q��<j��<6��<8��<:��<��<N��<���<'��<N��<^��<Y��<`   `   0��<4��<���<\��<*��<k��<B��<��<7��<:��<9��<<��<9��<0��<��<J��<f��<"��<a��<���<2��<,��<B��<B��<`   `   Z��<~��<K��<*��<���<N��<K��<>��<Z��<R��<P��<R��<a��<>��<?��<N��<���<*��<?��<~��<a��<'��<6��<'��<`   `   ���<U��<��<k��<N��<I��<J��<0��<c��<-��<*��<\��<0��<S��<M��<E��<f��<$��<Z��<~��<A��<c��<c��<C��<`   `   C��<E��<>��<B��<K��<J��<��<K��<G��< ��<P��<K��<���<J��<P��<B��<<��<E��<C��<F��<X��<���<V��<F��<`   `   ,��<o��<8��<��<>��<0��<K��<���<4��<.��<���<T��<0��<5��<��<?��<j��<'��<=��<X��<L��<O��<W��<8��<`   `   M��<8��<3��<7��<Z��<c��<G��<4��<9��<4��<A��<c��<c��<7��<(��<8��<V��<4��<j��<F��<@��<F��<p��<4��<`   `   G��<2��<j��<:��<R��<-��< ��<.��<4��<	��<*��<I��<9��<r��<6��<C��<Y��<L��<g��<���<���<b��<K��<_��<`   `   5��<^��<S��<9��<P��<*��<P��<���<A��<*��<\��<9��<M��<^��<5��<q��<V��<g��<k��<`��<s��<g��<Q��<q��<`   `   2��<g��<Q��<<��<R��<\��<K��<T��<c��<I��<9��<X��<g��<.��<?��<N��<V��<u��<T��<O��<r��<[��<M��<;��<`   `   j��<g��<Q��<9��<a��<0��<���<0��<c��<9��<M��<g��<o��<���<P��<C��<d��<[��<Y��<[��<a��<C��<T��<���<`   `   2��<a��<j��<0��<>��<S��<J��<5��<7��<r��<^��<.��<���<}��<6��<���<q��<H��<L��<v��<���<2��<}��<���<`   `   .��<6��<6��<��<?��<M��<P��<��<(��<6��<5��<?��<P��<6��<h��<^��<g��<���<]��<^��<o��<6��<P��<?��<`   `   G��<2��<8��<J��<N��<E��<B��<?��<8��<C��<q��<N��<C��<���<^��<��<k��<p��<��<Z��<���<C��<M��<t��<`   `   X��<j��<:��<f��<���<f��<<��<j��<V��<Y��<V��<V��<d��<q��<g��<k��<C��<k��<f��<q��<f��<V��<S��<Y��<`   `   ,��<M��<��<"��<*��<$��<E��<'��<4��<L��<g��<u��<[��<H��<���<p��<k��<���<L��<\��<r��<j��<K��<.��<`   `   6��<Z��<N��<a��<?��<Z��<C��<=��<j��<g��<k��<T��<Y��<L��<]��<��<f��<L��<T��<T��<k��<g��<q��<=��<`   `   ���<u��<���<���<~��<~��<F��<X��<F��<���<`��<O��<[��<v��<^��<Z��<q��<\��<T��<c��<���<@��<W��<N��<`   `   f��<2��<'��<2��<a��<A��<X��<L��<@��<���<s��<r��<a��<���<o��<���<f��<r��<k��<���<I��<L��<P��<A��<`   `   0��<U��<N��<,��<'��<c��<���<O��<F��<b��<g��<[��<C��<2��<6��<C��<V��<j��<g��<@��<L��<���<c��<��<`   `   S��<`��<^��<B��<6��<c��<V��<W��<p��<K��<Q��<M��<T��<}��<P��<M��<S��<K��<q��<W��<P��<c��<?��<B��<`   `   $��< ��<Y��<B��<'��<C��<F��<8��<4��<_��<q��<;��<���<���<?��<t��<Y��<.��<=��<N��<A��<��<B��<`��<`   `   ��<���<���<Շ�<���<���<���<Ň�<ڇ�<���<Շ�<���<���<���<Ӈ�<���<އ�<Ň�<���<���<���<Շ�<���<���<`   `   ���<f��<Ƈ�<���<V��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<Q��<���<ʇ�<d��<���<`   `   ���<Ƈ�<��<���<���<և�<���<���<͇�<���<���<ɇ�<���<���<Ӈ�<���<���<և�<���<���<އ�<Ƈ�<���<��<`   `   Շ�<���<���<���<���<�<Ç�<̇�<͇�<���<���<���<���<ȇ�<ˇ�<ȇ�<Ç�<���<���<���<���<ч�<݇�<߇�<`   `   ���<V��<���<���<���<���<���<ɇ�<���<���<χ�<���<���<ɇ�<���<���<���<���<���<V��<���<���<���<���<`   `   ���<���<և�<�<���<���<��<Ň�<���<݇�<ڇ�<���<Ǉ�<��<���<���<Ç�<ۇ�<���<���<Ň�<���<���<Ç�<`   `   ���<���<���<Ç�<���<��<���<���<���<���<���<���<���<��<���<Ç�<���<���<���<���<���<���<���<���<`   `   Ň�<���<���<̇�<ɇ�<Ň�<���<��<ʇ�<Ƈ�<���<���<Ǉ�<ć�<ˇ�<���<���<���<���<���<���<���<���<���<`   `   ڇ�<���<͇�<͇�<���<���<���<ʇ�<݇�<ʇ�<���<���<���<͇�<ʇ�<���<݇�<Ç�<���<���<���<���<���<Ç�<`   `   ���<���<���<���<���<݇�<���<Ƈ�<ʇ�<���<ڇ�<���<���<���<���<���<���<ć�<���<���<���<���<���<���<`   `   Շ�<���<���<���<χ�<ڇ�<���<���<���<ڇ�<ׇ�<���<���<���<ڇ�<���<���<���<q��<���<n��<���<���<���<`   `   ���<���<ɇ�<���<���<���<���<���<���<���<���<·�<���<���<ȇ�<���<���<h��<���<���<j��<���<���<ʇ�<`   `   ���<���<���<���<���<Ǉ�<���<Ǉ�<���<���<���<���<���<���<���<ڇ�<���<���<���<���<���<ڇ�<���<���<`   `   ���<���<���<ȇ�<ɇ�<��<��<ć�<͇�<���<���<���<���<���<���<���<���<���<���<���<���<���<~��<}��<`   `   Ӈ�<���<Ӈ�<ˇ�<���<���<���<ˇ�<ʇ�<���<ڇ�<ȇ�<���<���<s��<���<���<q��<���<���<p��<���<���<ȇ�<`   `   ���<���<���<ȇ�<���<���<Ç�<���<���<���<���<���<ڇ�<���<���<߇�<���<���<އ�<���<���<ׇ�<���<���<`   `   އ�<���<���<Ç�<���<Ç�<���<���<݇�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   Ň�<���<և�<���<���<ۇ�<���<���<Ç�<ć�<���<h��<���<���<q��<���<���<s��<���<���<j��<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<q��<���<���<���<���<އ�<���<���<���<���<l��<���<���<���<`   `   ���<Q��<���<���<V��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<އ�<���<���<Ň�<���<���<���<���<n��<j��<���<���<p��<���<���<j��<l��<���<���<���<���<Ň�<`   `   Շ�<ʇ�<Ƈ�<ч�<���<���<���<���<���<���<���<���<ڇ�<���<���<ׇ�<���<���<���<���<���<���<���<���<`   `   ���<d��<���<݇�<���<���<���<���<���<���<���<���<���<~��<���<���<���<���<���<���<���<���<���<݇�<`   `   ���<���<��<߇�<���<Ç�<���<���<Ç�<���<���<ʇ�<���<}��<ȇ�<���<���<���<���<���<Ň�<���<݇�<��<`   `   L��</��<��<)��<X��<��<!��<C��<.��<(��<:��<@��<r��<@��<=��<(��<)��<C��<'��<��<S��<)��<��</��<`   `   /��<D��<��<B��<6��<9��<��<���<#��<2��<��<��<��<��<,��<!��< ��<��<3��<5��<H��<��<?��<,��<`   `   ��<��<%��<��<3��<J��<��<A��<��<��<6��</��<.��<��<#��<A��<��<J��<;��<��<��<��<��<Ї�<`   `   )��<B��<��<(��<3��<��<@��<1��<��<B��</��<2��<F��<��<+��<A��<
��<2��<"��<��<H��<&��<���<��<`   `   X��<6��<3��<3��<��<B��<��<��<*��<��<��<��<'��<��<��<B��<���<3��<8��<6��<U��<<��<Z��<<��<`   `   ��<9��<J��<��<B��<+��<��<4��<��<<��<9��<��<9��<��<%��<A��<
��<K��<3��<��<��<O��<K��<��<`   `   !��<��<��<@��<��<��<]��<5��<��<>��<��<5��<W��<��<	��<@��<��<��<+��<!��<��<���<��<!��<`   `   C��<���<A��<1��<��<4��<5��<��<��< ��<��<6��<9��<��<+��<C��< ��<@��<9��<N��<X��<R��<J��<?��<`   `   .��<#��<��<��<*��<��<��<��<��<��<��<��<&��<��< ��<#��<*��<$��<��<6��<w��<6��<��<$��<`   `   (��<2��<��<B��<��<<��<>��< ��<��<?��<9��<��<F��<��<,��<%��<"��<3��< ��<#��<)��<��</��<��<`   `   :��<��<6��</��<��<9��<��<��<��<9��<��</��<0��<��<C��<&��<Q��<i��<`��<���<S��<i��<\��<&��<`   `   @��<��</��<2��<��<��<5��<6��<��<��</��<0��<��<>��<��<��<9��<O��<>��<E��<U��<2��<��<!��<`   `   r��<��<.��<F��<'��<9��<W��<9��<&��<F��<0��<��<p��<&��<��<��<?��<-��<��<-��<@��<��<��<&��<`   `   @��<��<��<��<��<��<��<��<��<��<��<>��<&��<Q��<c��<��<:��<K��<E��<3��<��<i��<L��<!��<`   `   =��<,��<#��<+��<��<%��<	��<+��< ��<,��<C��<��<��<c��<J��<Q��<:��<F��<G��<Q��<>��<c��<'��<��<`   `   (��<!��<A��<A��<B��<A��<@��<C��<#��<%��<&��<��<��<��<Q��<X��<-��<&��<Q��<W��<��<��<��<)��<`   `   )��< ��<��<
��<���<
��<��< ��<*��<"��<Q��<9��<?��<:��<:��<-��<L��<-��<:��<:��<>��<9��<R��<"��<`   `   C��<��<J��<2��<3��<K��<��<@��<$��<3��<i��<O��<-��<K��<F��<&��<-��<L��<E��<(��<U��<l��</��<"��<`   `   '��<3��<;��<"��<8��<3��<+��<9��<��< ��<`��<>��<��<E��<G��<Q��<:��<E��<��<>��<W��< ��<��<9��<`   `   ��<5��<��<��<6��<��<!��<N��<6��<#��<���<E��<-��<3��<Q��<W��<:��<(��<>��<���<)��<4��<J��<"��<`   `   S��<H��<��<H��<U��<��<��<X��<w��<)��<S��<U��<@��<��<>��<��<>��<U��<W��<)��<s��<X��<��<��<`   `   )��<��<��<&��<<��<O��<���<R��<6��<��<i��<2��<��<i��<c��<��<9��<l��< ��<4��<X��< ��<K��<;��<`   `   ��<?��<��<���<Z��<K��<��<J��<��</��<\��<��<��<L��<'��<��<R��</��<��<J��<��<K��<_��<���<`   `   /��<,��<Ї�<��<<��<��<!��<?��<$��<��<&��<!��<&��<!��<��<)��<"��<"��<9��<"��<��<;��<���<҇�<`   `   ��<���<��<���<���<���<���<���<���<���<���<���<ʈ�<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<��<���<���<ۈ�<���<���<���<���<҈�<È�<���<���<ň�<Ȉ�<���<���<���<���<߈�<���<���<
��<���<`   `   ��<���<���<ň�<���<���<ވ�<���<���<���<ψ�<���<ň�<���<���<���<Ո�<���<���<ň�<���<���<���<���<`   `   ���<���<ň�<���<È�<���<���<ň�<���<È�<���<���<ʈ�<���<���<���<���<ǈ�<���<È�<���<���<߈�<��<`   `   ���<ۈ�<���<È�<܈�<ǈ�<���<��<݈�<���<���<���<Ո�<��<Ɉ�<ǈ�<͈�<È�<���<ۈ�<���<p��<���<p��<`   `   ���<���<���<���<ǈ�<���<���<���<���<���<���<���<���<���<��<ˈ�<���<���<���<���<���<ƈ�<���<���<`   `   ���<���<ވ�<���<���<���<���<���<���<���<���<���<���<���<�<���<Ԉ�<���<���<���<���<���<���<���<`   `   ���<���<���<ň�<��<���<���<߈�<ш�<҈�<܈�<���<���<��<���<���<���<���<���<���<���<|��<���<Ȉ�<`   `   ���<���<���<���<݈�<���<���<ш�<��<ш�<���<���<҈�<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<҈�<���<È�<���<���<���<҈�<ш�<���<���<Ĉ�<ʈ�<���<Ȉ�<���<���<���<Ȉ�<t��<}��<ӈ�<���<���<`   `   ���<È�<ψ�<���<���<���<���<܈�<���<���<���<���<ʈ�<È�<���<���<���<t��<���<���<���<t��<���<���<`   `   ���<���<���<���<���<���<���<���<���<Ĉ�<���<���<���<���<���<҈�<x��<���<���<���<���<l��<͈�<���<`   `   ʈ�<���<ň�<ʈ�<Ո�<���<���<���<҈�<ʈ�<ʈ�<���<ň�<���<���<���<ۈ�<���<T��<���<ވ�<���<���<���<`   `   ���<ň�<���<���<��<���<���<��<���<���<È�<���<���<���<���<���<���<ӈ�<Ȉ�<���<���<���<���<���<`   `   ���<Ȉ�<���<���<Ɉ�<��<�<���<���<Ȉ�<���<���<���<���<���<���<l��<ˈ�<���<���<���<���<���<���<`   `   ���<���<���<���<ǈ�<ˈ�<���<���<���<���<���<҈�<���<���<���<b��<���<���<V��<���<���<���<͈�<���<`   `   ���<���<Ո�<���<͈�<���<Ԉ�<���<���<���<���<x��<ۈ�<���<l��<���<��<���<n��<���<و�<x��<���<���<`   `   ���<���<���<ǈ�<È�<���<���<���<���<���<t��<���<���<ӈ�<ˈ�<���<���<Ո�<Ȉ�<���<���<v��<���<���<`   `   ���<���<���<���<���<���<���<���<���<Ȉ�<���<���<T��<Ȉ�<���<V��<n��<Ȉ�<f��<���<���<Ȉ�<���<���<`   `   ���<߈�<ň�<È�<ۈ�<���<���<���<���<t��<���<���<���<���<���<���<���<���<���<���<}��<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<}��<���<���<ވ�<���<���<���<و�<���<���<}��<���<���<���<���<`   `   ���<���<���<���<p��<ƈ�<���<|��<���<ӈ�<t��<l��<���<���<���<���<x��<v��<Ȉ�<���<���<���<���<s��<`   `   ���<
��<���<߈�<���<���<���<���<���<���<���<͈�<���<���<���<͈�<���<���<���<���<���<���<���<߈�<`   `   ���<���<���<��<p��<���<���<Ȉ�<���<���<���<���<���<���<���<���<���<���<���<���<���<s��<߈�<���<`   `   	��<O��<��<m��<[��<U��<C��<C��<q��<V��<)��<Q��<M��<Q��<5��<V��<]��<C��<Z��<U��<G��<m��<��<O��<`   `   O��<��<Q��<3��<1��<l��<Y��<)��<G��<v��<f��<T��<\��<h��<i��<K��<9��<P��<]��<9��<>��<K��<	��<P��<`   `   ��<Q��<���<F��<)��<Z��<���<?��<:��<D��<I��<J��<@��<D��<C��<?��<���<Z��</��<F��<���<Q��<��<���<`   `   m��<3��<F��<b��<V��<5��<*��<o��<L��<���<M��<N��<��<P��<b��<"��<E��<_��<R��<@��<>��<n��<a��<g��<`   `   [��<1��<)��<V��<o��<!��<��<b��<��<I��<k��<I��<��<b��<&��<!��<W��<V��<>��<1��<O��<l��<
��<l��<`   `   U��<l��<Z��<5��<!��<*��<V��<,��<H��<S��<R��<M��<4��<N��<��<*��<E��<T��<]��<V��<s��<H��<B��<h��<`   `   C��<Y��<���<*��<��<V��<q��<I��<S��<#��<P��<I��<r��<V��<��<*��<���<Y��<Q��<R��<e��<m��<v��<R��<`   `   C��<)��<?��<o��<b��<,��<I��<P��<*��<.��<O��<A��<4��<k��<b��<9��<9��<D��<E��<#��<F��<;��<��<T��<`   `   q��<G��<:��<L��<��<H��<S��<*��<��<*��<]��<H��<	��<L��<N��<G��<a��<S��<6��<o��<���<o��<,��<S��<`   `   V��<v��<D��<���<I��<S��<#��<.��<*��<��<R��<R��<��<>��<i��<W��<F��<U��<���<U��<`��<���<O��<6��<`   `   )��<f��<I��<M��<k��<R��<P��<O��<]��<R��<c��<M��<H��<f��<5��<?��<<��<J��<a��<T��<F��<J��<R��<?��<`   `   Q��<T��<J��<N��<I��<M��<I��<A��<H��<R��<M��<C��<\��<R��<o��<u��<Z��<E��<���<���<P��<K��<p��<|��<`   `   M��<\��<@��<��<��<4��<r��<4��<	��<��<H��<\��<D��<@��<W��<e��<���<S��<q��<S��<���<e��<O��<@��<`   `   Q��<h��<D��<P��<b��<N��<V��<k��<L��<>��<f��<R��<@��<I��<]��<K��<��<Z��<K��<��<W��<j��<D��<8��<`   `   5��<i��<C��<b��<&��<��<��<b��<N��<i��<5��<o��<W��<]��<���<���<?��<Q��<^��<���<j��<]��<d��<o��<`   `   V��<K��<?��<"��<!��<*��<*��<9��<G��<W��<?��<u��<e��<K��<���<؉�<[��<K��<ɉ�<���<W��<^��<p��<A��<`   `   ]��<9��<���<E��<W��<E��<���<9��<a��<F��<<��<Z��<���<��<?��<[��<\��<[��<A��<��<���<Z��<A��<F��<`   `   C��<P��<Z��<_��<V��<T��<Y��<D��<S��<U��<J��<E��<S��<Z��<Q��<K��<[��<^��<K��<K��<P��<K��<O��<W��<`   `   Z��<]��</��<R��<>��<]��<Q��<E��<6��<���<a��<���<q��<K��<^��<ɉ�<A��<K��<���<���<T��<���<7��<E��<`   `   U��<9��<F��<@��<1��<V��<R��<#��<o��<U��<T��<���<S��<��<���<���<��<K��<���<V��<`��<s��<��<I��<`   `   G��<>��<���<>��<O��<s��<e��<F��<���<`��<F��<P��<���<W��<j��<W��<���<P��<T��<`��<u��<F��<s��<s��<`   `   m��<K��<Q��<n��<l��<H��<m��<;��<o��<���<J��<K��<e��<j��<]��<^��<Z��<K��<���<s��<F��<e��<B��<u��<`   `   ��<	��<��<a��<
��<B��<v��<��<,��<O��<R��<p��<O��<D��<d��<p��<A��<O��<7��<��<s��<B��<��<a��<`   `   O��<P��<���<g��<l��<h��<R��<T��<S��<6��<?��<|��<@��<8��<o��<A��<F��<W��<E��<I��<s��<u��<a��<��<`   `   ���<���<���<��<��<ۉ�<݉�<���<*��<���<Չ�<��<���<��<��<���<��<���<���<ۉ�<׉�<��<��<���<`   `   ���<��< ��<���<��<I��<ĉ�<���<���<���<ى�<��<��<ى�<��<��<ʉ�<���<7��<��<ǉ�<��<��<��<`   `   ���< ��<!��<��<��<̉�<��<��<��<���<	��<	��<��<���<��<��<��<̉�<��<��<��< ��<���<���<`   `   ��<���<��<9��<܉�<щ�<(��<��<(��<!��<��<��<)��<0��<��<��<��<��<'��<ى�<ǉ�<
��<��<��<`   `   ��<��<��<܉�<
��<Q��<��<މ�<��<$��<���<$��<��<މ�<��<Q��<��<܉�<*��<��<��<,��<щ�<,��<`   `   ۉ�<I��<̉�<щ�<Q��</��<��<���<%��<ى�<ى�<-��<��<��<!��<_��<��<�<7��<߉�<ى�<��<��<͉�<`   `   ݉�<ĉ�<��<(��<��<��<F��<��<��<"��<��<��<K��<��<��<(��<��<ĉ�<��<؉�<��<��<��<؉�<`   `   ���<���<��<��<މ�<���<��<ŉ�<&��<.��<ŉ�<���<��<��<��<݉�<ʉ�<���<?��<��<���<���<��<P��<`   `   *��<���<��<(��<��<%��<��<&��<��<&��< ��<%��<���<(��<���<���<��<��<���<��<��<��<���<��<`   `   ���<���<���<!��<$��<ى�<"��<.��<&��<��<ى�<1��<)��<��<��<��<��<��<ω�<�<Ή�<���<܉�<ډ�<`   `   Չ�<ى�<	��<��<���<ى�<��<ŉ�< ��<ى�<���<��<��<ى�<��<��<��<(��<��<��<Љ�<(��</��<��<`   `   ��<��<	��<��<$��<-��<��<���<%��<1��<��<���<��<��<��<���<���<ω�<݉�<��<ۉ�<��<���<%��<`   `   ���<��<��<)��<��<��<K��<��<���<)��<��<��<���<���<���<���<!��<���<���<���<&��<���<���<���<`   `   ��<ى�<���<0��<މ�<��<��<��<(��<��<ى�<��<���<��<��<݉�<��<,��<��<���<��<'��<��<���<`   `   ��<��<��<��<��<!��<��<��<���<��<��<��<���<��<�<���<��<���<��<���<���<��<ĉ�<��<`   `   ���<��<��<��<Q��<_��<(��<݉�<���<��<��<���<���<݉�<���<��<Ή�<���<��<É�<��<���<���<��<`   `   ��<ʉ�<��<��<��<��<��<ʉ�<��<��<��<���<!��<��<��<Ή�<���<Ή�<��<��<��<���<��<��<`   `   ���<���<̉�<��<܉�<�<ĉ�<���<��<��<(��<ω�<���<,��<���<���<Ή�<��<��<���<ۉ�<(��<܉�<��<`   `   ���<7��<��<'��<*��<7��<��<?��<���<ω�<��<݉�<���<��<��<��<��<��<؉�<݉�<��<ω�<���<?��<`   `   ۉ�<��<��<ى�<��<߉�<؉�<��<��<�<��<��<���<���<���<É�<��<���<݉�<��<Ή�<��<��<ˉ�<`   `   ׉�<ǉ�<��<ǉ�<��<ى�<��<���<��<Ή�<Љ�<ۉ�<&��<��<���<��<��<ۉ�<��<Ή�<��<���<��<ى�<`   `   ��<��< ��<
��<,��<��<��<���<��<���<(��<��<���<'��<��<���<���<(��<ω�<��<���<׉�<��<:��<`   `   ��<��<���<��<щ�<��<��<��<���<܉�</��<���<���<��<ĉ�<���<��<܉�<���<��<��<��<ȉ�<��<`   `   ���<��<���<��<,��<͉�<؉�<P��<��<ډ�<��<%��<���<���<��<��<��<��<?��<ˉ�<ى�<:��<��<��<`   `   ى�<���<Ȋ�<���<܊�<���<���<���<Ê�<���<���<���<���<���<���<���<���<���<���<���<���<���<ي�<���<`   `   ���<ϊ�<���<���<��<ڊ�<ϊ�<Њ�<��<���<Ċ�<���<���<�<���<���<��<���<Ǌ�<���<���<v��<ˊ�<Ɗ�<`   `   Ȋ�<���<��<���<q��<���<'��<���<���<���<Ŋ�<���<���<���<���<���<$��<���<r��<���<���<���<Ɗ�<��<`   `   ���<���<���<׊�<��<���<���<���<���<���<���<���<���<���<���<���<���<���<Ŋ�<���<���<���<���<���<`   `   ܊�<��<q��<��<���<���<���<ي�<���<̊�<���<̊�<���<ي�<���<���<���<��<���<��<Ɋ�<Ǌ�<���<Ǌ�<`   `   ���<ڊ�<���<���<���<���<���<���<���<���<���<Ê�<���<���<���<���<���<���<Ǌ�<Ǌ�<���<��<��<���<`   `   ���<ϊ�<'��<���<���<���<��<���<���<���<���<���<��<���<���<���<!��<ϊ�<���<���<؊�<���<��<���<`   `   ���<Њ�<���<���<ي�<���<���<���<���<���<���<���<���<��<���<���<��<���<Ҋ�<��<���<���<��<��<`   `   Ê�<��<���<���<���<���<���<���<T��<���<ʊ�<���<���<���<���<��<���<���<���<ъ�<ϊ�<ъ�<���<���<`   `   ���<���<���<���<̊�<���<���<���<���<���<���<ފ�<���<���<���<���<���<Ɋ�<��<Ȋ�<Պ�<���<Ŋ�<���<`   `   ���<Ċ�<Ŋ�<���<���<���<���<���<ʊ�<���<���<���<̊�<Ċ�<���<ϊ�<Њ�<���<ߊ�<��<���<���<��<ϊ�<`   `   ���<���<���<���<̊�<Ê�<���<���<���<ފ�<���<���<���<���<��<��<���<���<���<	��<���<���<���<���<`   `   ���<���<���<���<���<���<��<���<���<���<̊�<���<���<���<���<ˊ�<���<���<���<���<��<ˊ�<���<���<`   `   ���<�<���<���<ي�<���<���<��<���<���<Ċ�<���<���<�<ي�<׊�<��<���<͊�<ڊ�<��<��<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<��<���<ي�<���<��<���<���<͊�<��<���<ي�<Ɗ�<��<`   `   ���<���<���<���<���<���<���<���<��<���<ϊ�<��<ˊ�<׊�<��<Պ�<Ċ�<���<�<���<��<Ċ�<���<͊�<`   `   ���<��<$��<���<���<���<!��<��<���<���<Њ�<���<���<��<���<Ċ�<���<Ċ�<���<��<���<���<׊�<���<`   `   ���<���<���<���<��<���<ϊ�<���<���<Ɋ�<���<���<���<���<���<���<Ċ�<���<͊�<���<���<���<Ŋ�<���<`   `   ���<Ǌ�<r��<Ŋ�<���<Ǌ�<���<Ҋ�<���<��<ߊ�<���<���<͊�<͊�<�<���<͊�<���<���<Ԋ�<��<���<Ҋ�<`   `   ���<���<���<���<��<Ǌ�<���<��<ъ�<Ȋ�<��<	��<���<ڊ�<��<���<��<���<���<��<Պ�<݊�<��<���<`   `   ���<���<���<���<Ɋ�<���<؊�<���<ϊ�<Պ�<���<���<��<��<���<��<���<���<Ԋ�<Պ�<���<���<��<���<`   `   ���<v��<���<���<Ǌ�<��<���<���<ъ�<���<���<���<ˊ�<��<ي�<Ċ�<���<���<��<݊�<���<���<��<؊�<`   `   ڊ�<ˊ�<Ɗ�<���<���<��<��<��<���<Ŋ�<��<���<���<���<Ɗ�<���<׊�<Ŋ�<���<��<��<��<���<���<`   `   ���<Ɗ�<��<���<Ǌ�<���<���<��<���<���<ϊ�<���<���<���<��<͊�<���<���<Ҋ�<���<���<؊�<���<��<`   `   ��<���<p��<���<���<���<���<���<���<���<I��<���<Ë�<���<\��<���<s��<���<���<���<j��<���<���<���<`   `   ���<���<���<���<���<���<��<@��<���<���<���<���<���<���<���<���<S��<k��<���<���<���<p��<���<���<`   `   p��<���<��<���<7��<~��<Ë�<Z��<y��<���<ŋ�<���<Ë�<���<z��<Z��<ċ�<~��<5��<���<��<���<j��<6��<`   `   ���<���<���<���<���<}��<t��<ċ�<���<l��<���<���<s��<���<���<`��<���<Ӌ�<���<v��<���<Ë�<���<���<`   `   ���<���<7��<���<���<���<���<Ћ�<v��<���<�<���<a��<Ћ�<���<���<~��<���<Z��<���<w��<���<���<���<`   `   ���<���<~��<}��<���<Ƌ�<l��<���<���<���<���<���<���<X��<���<͋�<���<n��<���<���<j��<n��<k��<^��<`   `   ���<��<Ë�<t��<���<l��<���<���<���<g��<���<���<���<l��<���<t��<���<��<���<���<���<z��<���<���<`   `   ���<@��<Z��<ċ�<Ћ�<���<���<���<���<���<ŋ�<���<���<��<���<J��<S��<���<p��<d��<���<���<a��<���<`   `   ���<���<y��<���<v��<���<���<���<p��<���<���<���<Z��<���<���<���<y��<���<P��<���<���<���<@��<���<`   `   ���<���<���<l��<���<���<g��<���<���<S��<���<���<s��<w��<���<���<���<���<���<Y��<e��<���<���<���<`   `   I��<���<ŋ�<���<�<���<���<ŋ�<���<���<���<���<ϋ�<���<P��<{��<x��<c��<z��<��<Z��<c��<���<{��<`   `   ���<���<���<���<���<���<���<���<���<���<���<t��<���<���<q��<���<p��<���<���<���<���<\��<���<���<`   `   Ë�<���<Ë�<s��<a��<���<���<���<Z��<s��<ϋ�<���<���<���<~��<���<���<���<V��<���<���<���<q��<���<`   `   ���<���<���<���<Ћ�<X��<l��<��<���<w��<���<���<���<���<v��<*��< ��<���<���<��<6��<���<���<���<`   `   \��<���<z��<���<���<���<���<���<���<���<P��<q��<~��<v��<v��<���<f��<���<���<���<[��<v��<���<q��<`   `   ���<���<Z��<`��<���<͋�<t��<J��<���<���<{��<���<���<*��<���<���<N��<:��<���<�<6��<���<���<w��<`   `   s��<S��<ċ�<���<~��<���<���<S��<y��<���<x��<p��<���< ��<f��<N��<���<N��<j��< ��<���<p��<��<���<`   `   ���<k��<~��<Ӌ�<���<n��<��<���<���<���<c��<���<���<���<���<:��<N��<Ë�<���<z��<���<^��<���<���<`   `   ���<���<5��<���<Z��<���<���<p��<P��<���<z��<���<V��<���<���<���<j��<���<o��<���<q��<���<E��<p��<`   `   ���<���<���<v��<���<���<���<d��<���<Y��<��<���<���<��<���<�< ��<z��<���<��<e��<���<a��<v��<`   `   j��<���<��<���<w��<j��<���<���<���<e��<Z��<���<���<6��<[��<6��<���<���<q��<e��<���<���<ɋ�<j��<`   `   ���<p��<���<Ë�<���<n��<z��<���<���<���<c��<\��<���<���<v��<���<p��<^��<���<���<���<f��<k��<���<`   `   ���<���<j��<���<���<k��<���<a��<@��<���<���<���<q��<���<���<���<��<���<E��<a��<ɋ�<k��<u��<���<`   `   ���<���<6��<���<���<^��<���<���<���<���<{��<���<���<���<q��<w��<���<���<p��<v��<j��<���<���<%��<`   `   Z��<W��<���<���<5��<��<[��<���<���<���<���<���<}��<���<���<���<j��<���<���<��<��<���<���<W��<`   `   W��<���<i��<��<���<���<@��<O��<���<r��<Y��<+��<0��<S��<d��<���<a��<*��<���<���<"��<V��<���<a��<`   `   ���<i��<V��<i��<���<w��<���<���<i��<?��<���<K��<���<?��<h��<���<���<w��<���<i��<]��<i��<���<1��<`   `   ���<��<i��<���<D��<F��<d��<���<t��<���<W��<Q��<���<���<s��<N��<X��<[��<���<W��<"��<���<���<���<`   `   5��<���<���<D��<��<���<��<F��<r��<y��<��<y��<]��<F��<:��<���<��<D��<���<���< ��<���<n��<���<`   `   ��<���<w��<F��<���<���<E��<}��<���<a��<g��<���<���</��<���<���<X��<d��<���<���<^��<g��<f��<R��<`   `   [��<@��<���<d��<��<E��<Ì�<?��<l��<j��<V��<?��<Ԍ�<E��<��<d��<���<@��<c��<s��<���<S��<���<s��<`   `   ���<O��<���<���<F��<}��<?��<5��<x��<���<:��<)��<���<]��<s��<��<a��<���<���<���<n��<c��<���<���<`   `   ���<���<i��<t��<r��<���<l��<x��<)��<x��<|��<���<V��<t��<���<���<p��<���<H��<{��<���<{��<8��<���<`   `   ���<r��<?��<���<y��<a��<j��<���<x��<T��<g��<���<���<-��<d��<���<O��<k��<���<���<���<���<j��<<��<`   `   ���<Y��<���<W��<��<g��<V��<:��<|��<g��<���<W��<���<Y��<���<���<���<l��<���<���<��<l��<���<���<`   `   ���<+��<K��<Q��<y��<���<?��<)��<���<���<W��<8��<0��<���<x��<o��<j��<}��<z��<���<���<W��<n��<���<`   `   }��<0��<���<���<]��<���<Ԍ�<���<V��<���<���<0��<o��<v��<L��<���<Č�<���<#��<���<̌�<���<@��<v��<`   `   ���<S��<?��<���<F��</��<E��<]��<t��<-��<Y��<���<v��<���<���<s��<v��<���<���<d��<~��<���<���<q��<`   `   ���<d��<h��<s��<:��<���<��<s��<���<d��<���<x��<L��<���<���<���<d��<�<���<���<���<���<S��<x��<`   `   ���<���<���<N��<���<���<d��<��<���<���<���<o��<���<s��<���<u��<t��<a��<c��<���<~��<���<n��<���<`   `   j��<a��<���<X��<��<X��<���<a��<p��<O��<���<j��<Č�<v��<d��<t��<��<t��<h��<v��<���<j��<���<O��<`   `   ���<*��<w��<[��<D��<d��<@��<���<���<k��<l��<}��<���<���<�<a��<t��<Ќ�<���<���<���<f��<j��<���<`   `   ���<���<���<���<���<���<c��<���<H��<���<���<z��<#��<���<���<c��<h��<���<:��<z��<���<���<:��<���<`   `   ��<���<i��<W��<���<���<s��<���<{��<���<���<���<���<d��<���<���<v��<���<z��<���<���<���<���<]��<`   `   ��<"��<]��<"��< ��<^��<���<n��<���<���<��<���<̌�<~��<���<~��<���<���<���<���<i��<n��<Ì�<^��<`   `   ���<V��<i��<���<���<g��<S��<c��<{��<���<l��<W��<���<���<���<���<j��<f��<���<���<n��<=��<f��<���<`   `   ���<���<���<���<n��<f��<���<���<8��<j��<���<n��<@��<���<S��<n��<���<j��<:��<���<Ì�<f��<Y��<���<`   `   W��<a��<1��<���<���<R��<s��<���<���<<��<���<���<v��<q��<x��<���<O��<���<���<]��<^��<���<���<��<`   `   :��<��<y��<L��<���<���<!��<���<U��<Z��<V��<y��<l��<y��<i��<Z��<4��<���<G��<���<o��<L��<���<��<`   `   ��<C��<]��<x��<���<b��<F��<K��<m��<o��<o��<��<���<h��<c��<}��<\��</��<R��<���<���<J��<C��<���<`   `   y��<]��<ߍ�<\��< ��<b��<���<F��<S��<D��<���<|��<���<D��<N��<F��<���<b��<��<\��<��<]��<n��<���<`   `   L��<x��<\��<`��<���<w��<B��<���<���<U��<r��<k��<Y��<���<���<+��<���<���<Q��<I��<���<V��<*��<*��<`   `   ���<���< ��<���<���<w��<Q��<���<6��<|��<���<|��<"��<���<t��<w��<f��<���<B��<���<|��<k��<(��<k��<`   `   ���<b��<b��<w��<w��<���<���<b��<v��<}��<���<���<f��<o��<���<���<���<O��<R��<���<���<���<���<{��<`   `   !��<F��<���<B��<Q��<���<���<I��<���<V��<}��<I��<���<���<F��<B��<���<F��<&��<��<l��<5��<v��<��<`   `   ���<K��<F��<���<���<b��<I��<���<���<���<���<2��<f��<���<���<3��<\��<���<l��<���<M��<C��<���<|��<`   `   U��<m��<S��<���<6��<v��<���<���<��<���<���<v��<��<���<r��<m��<:��<N��<Z��<}��<P��<}��<J��<N��<`   `   Z��<o��<D��<U��<|��<}��<V��<���<���<?��<���<���<Y��<1��<c��<d��<��<t��<`��<5��<?��<p��<t��<	��<`   `   V��<o��<���<r��<���<���<}��<���<���<���<h��<r��<���<o��<W��<W��<���<s��<V��<���<<��<s��<ō�<W��<`   `   y��<��<|��<k��<|��<���<I��<2��<v��<���<r��<i��<���<���<f��<l��<8��< ��<w��<���<
��<'��<l��<r��<`   `   l��<���<���<Y��<"��<f��<���<f��<��<Y��<���<���<^��<T��<_��<O��<i��<a��<;��<a��<p��<O��<S��<T��<`   `   y��<h��<D��<���<���<o��<���<���<���<1��<o��<���<T��<_��<V��<C��<u��<[��<K��<e��<L��<b��<_��<P��<`   `   i��<c��<N��<���<t��<���<F��<���<r��<c��<W��<f��<_��<V��<��<f��</��<��<O��<f��<��<V��<c��<f��<`   `   Z��<}��<F��<+��<w��<���<B��<3��<m��<d��<W��<l��<O��<C��<f��<���<M��<<��<���<s��<L��<K��<l��<P��<`   `   4��<\��<���<���<f��<���<���<\��<:��<��<���<8��<i��<u��</��<M��<���<M��<2��<u��<c��<8��<���<��<`   `   ���</��<b��<���<���<O��<F��<���<N��<t��<s��< ��<a��<[��<��<<��<M��<��<K��<]��<
��<l��<t��<^��<`   `   G��<R��<��<Q��<B��<R��<&��<l��<Z��<`��<V��<w��<;��<K��<O��<���<2��<K��<N��<w��<S��<`��<J��<l��<`   `   ���<���<\��<I��<���<���<��<���<}��<5��<���<���<a��<e��<f��<s��<u��<]��<w��<���<?��<���<���<���<`   `   o��<���<��<���<|��<���<l��<M��<P��<?��<<��<
��<p��<L��<��<L��<c��<
��<S��<?��<7��<M��<���<���<`   `   L��<J��<]��<V��<k��<���<5��<C��<}��<p��<s��<'��<O��<b��<V��<K��<8��<l��<`��<���<M��<��<���<���<`   `   ���<C��<n��<*��<(��<���<v��<���<J��<t��<ō�<l��<S��<_��<c��<l��<���<t��<J��<���<���<���<��<*��<`   `   ��<���<���<*��<k��<{��<��<|��<N��<	��<W��<r��<T��<P��<f��<P��<��<^��<l��<���<���<���<*��<���<`   `   P��<r��<{��<|��<P��<���<���<���<���<���<8��<b��<l��<b��<I��<���<���<���<���<���<3��<|��<���<r��<`   `   r��<S��<V��<N��<a��<���<���<M��<���<���<e��<e��<g��<^��<���<���<[��<u��<���<w��<U��<D��<T��<}��<`   `   {��<V��<���<O��<2��<Q��<���<9��<W��<~��<j��<��<o��<~��<R��<9��<���<Q��<)��<O��<���<V��<p��<r��<`   `   |��<N��<O��<���<���<2��<`��<���<���<[��<W��<P��<]��<���<���<K��<@��<���<���<=��<U��<���<���<���<`   `   P��<a��<2��<���<D��<m��<s��<���<H��<���<���<���<6��<���<���<m��< ��<���<Q��<a��<>��<���<~��<���<`   `   ���<���<Q��<2��<m��<p��<*��<`��<���<>��<E��<���<c��<��<f��<���<@��<?��<���<���<M��<j��<k��<F��<`   `   ���<���<���<`��<s��<*��<h��<g��<q��<��<Z��<g��<z��<*��<g��<`��<���<���<���<\��<s��<Z��<z��<\��<`   `   ���<M��<9��<���<���<`��<g��<v��<���<���<}��<R��<c��<���<���<'��<[��<���<���<���<���<���<���<���<`   `   ���<���<W��<���<H��<���<q��<���<M��<���<��<���<0��<���<s��<���<���<���<J��<���<���<���<<��<���<`   `   ���<���<~��<[��<���<>��<��<���<���<���<E��<���<]��<l��<���<Î�<���<}��<h��<_��<g��<u��<~��<���<`   `   8��<e��<j��<W��<���<E��<Z��<}��<��<E��<~��<W��<z��<e��<8��<H��<���<���<���<`��<l��<���<���<H��<`   `   b��<e��<��<P��<���<���<g��<R��<���<���<W��<	��<g��<m��<��<f��<n��<���<���<���<���<`��<g��<���<`   `   l��<g��<o��<]��<6��<c��<z��<c��<0��<]��<z��<g��<_��<|��<���<���<���<���<p��<���<���<���<���<|��<`   `   b��<^��<~��<���<���<��<*��<���<���<l��<e��<m��<|��<s��<���<z��<S��<���<���<E��<���<���<t��<z��<`   `   I��<���<R��<���<���<f��<g��<���<s��<���<8��<��<���<���<���<���<t��<ǎ�<���<���<��<���<���<��<`   `   ���<���<9��<K��<m��<���<`��<'��<���<Î�<H��<f��<���<z��<���<���<y��<k��<���<���<���<���<g��<A��<`   `   ���<[��<���<@��< ��<@��<���<[��<���<���<���<n��<���<S��<t��<y��<J��<y��<w��<S��<���<n��<���<���<`   `   ���<u��<Q��<���<���<?��<���<���<���<}��<���<���<���<���<ǎ�<k��<y��<ю�<���<���<���<���<~��<���<`   `   ���<���<)��<���<Q��<���<���<���<J��<h��<���<���<p��<���<���<���<w��<���<���<���<���<h��<:��<���<`   `   ���<w��<O��<=��<a��<���<\��<���<���<_��<`��<���<���<E��<���<���<S��<���<���<Y��<g��<���<���<G��<`   `   3��<U��<���<U��<>��<M��<s��<���<���<g��<l��<���<���<���<��<���<���<���<���<g��<���<���<���<M��<`   `   |��<D��<V��<���<���<j��<Z��<���<���<u��<���<`��<���<���<���<���<n��<���<h��<���<���<E��<k��<���<`   `   ���<T��<p��<���<~��<k��<z��<���<<��<~��<���<g��<���<t��<���<g��<���<~��<:��<���<���<k��<g��<���<`   `   r��<}��<r��<���<���<F��<\��<���<���<���<H��<���<|��<z��<��<A��<���<���<���<G��<M��<���<���<`��<`   `   ���<���<���<���<m��<���<`��<>��<b��<~��<x��<���<���<���<���<~��<J��<>��<|��<���<U��<���<���<���<`   `   ���<֏�<���<~��<���<���<V��<p��<���<���<���<���<���<{��<}��<���<{��<D��<���<̏�<���<w��<؏�<���<`   `   ���<���<���<���<���<p��<���<���<l��<���<���<���<���<���<f��<���<���<p��<���<���<���<���<���<��<`   `   ���<~��<���<Ǐ�<���<b��<���<o��<}��<���<���<���<���<���<g��<���<m��<���<���<���<���<Ï�<���<���<`   `   m��<���<���<���<���<Џ�<r��<~��<{��<���<q��<���<l��<~��<���<Џ�<e��<���<ɏ�<���<^��<���<b��<���<`   `   ���<���<p��<b��<Џ�<���<���<���<���<���<���<���<���<{��<���<��<m��<`��<���<���<���<u��<w��<���<`   `   `��<V��<���<���<r��<���<���<���<���<��<���<���<��<���<g��<���<���<V��<a��<���<Ϗ�<���<ԏ�<���<`   `   >��<p��<���<o��<~��<���<���<+��<���<���<2��<m��<���<���<g��<���<{��<G��<���<p��<V��<Q��<r��<���<`   `   b��<���<l��<}��<{��<���<���<���<Q��<���<���<���<g��<}��<���<���<N��<���<u��<{��<f��<{��<i��<���<`   `   ~��<���<���<���<���<���<��<���<���<Џ�<���<���<���<z��<}��<���<���<p��<���<���<���<���<q��<��<`   `   x��<���<���<���<q��<���<���<2��<���<���<X��<���<Ï�<���<w��<���<i��<b��<���<���<���<b��<r��<���<`   `   ���<���<���<���<���<���<���<m��<���<���<���<���<���<���<͏�<���<p��<���<r��<|��<���<e��<���<Տ�<`   `   ���<���<���<���<l��<���<��<���<g��<���<Ï�<���<~��<x��<r��<c��<���<l��<H��<l��<���<c��<i��<x��<`   `   ���<{��<���<���<~��<{��<���<���<}��<z��<���<���<x��<J��<s��<���<R��<���<}��<G��<���<{��<K��<w��<`   `   ���<}��<f��<g��<���<���<g��<g��<���<}��<w��<͏�<r��<s��<���<y��<L��<���<b��<y��<���<s��<r��<͏�<`   `   ~��<���<���<���<Џ�<��<���<���<���<���<���<���<c��<���<y��<i��<}��<r��<_��<���<���<b��<���<���<`   `   J��<{��<���<m��<e��<m��<���<{��<N��<���<i��<p��<���<R��<L��<}��<���<}��<O��<R��<���<p��<n��<���<`   `   >��<D��<p��<���<���<`��<V��<G��<���<p��<b��<���<l��<���<���<r��<}��<���<}��<j��<���<\��<q��<���<`   `   |��<���<���<���<ɏ�<���<a��<���<u��<���<���<r��<H��<}��<b��<_��<O��<}��<S��<r��<���<���<f��<���<`   `   ���<̏�<���<���<���<���<���<p��<{��<���<���<|��<l��<G��<y��<���<R��<j��<r��<z��<���<���<r��<���<`   `   U��<���<���<���<^��<���<Ϗ�<V��<f��<���<���<���<���<���<���<���<���<���<���<���<S��<V��<���<���<`   `   ���<w��<���<Ï�<���<u��<���<Q��<{��<���<b��<e��<c��<{��<s��<b��<p��<\��<���<���<V��<���<w��<���<`   `   ���<؏�<���<���<b��<w��<ԏ�<r��<i��<q��<r��<���<i��<K��<r��<���<n��<q��<f��<r��<���<w��<N��<���<`   `   ���<���<��<���<���<���<���<���<���<��<���<Տ�<x��<w��<͏�<���<���<���<���<���<���<���<���<��<`   `   r��<֐�<���<���<���<���<���<
��<А�<���<���<���<���<���<���<���<���<
��<Ԑ�<���<���<���<���<֐�<`   `   ֐�<���<���<ؐ�<̐�<���<���<ϐ�<Ӑ�<ߐ�<���<���<���<���<ِ�<ސ�<א�<���<���<ڐ�<ܐ�<}��<���<ݐ�<`   `   ���<���<���<���<���<���<�<���<А�<���<���<���<���<���<ː�<���<Ȑ�<���<���<���<���<���<���<��<`   `   ���<ؐ�<���<W��<Ր�<���<o��<֐�<��<���<���<���<���<��<ѐ�<b��<���<��<P��<~��<ܐ�<���<͐�<ː�<`   `   ���<̐�<���<Ր�<���<���<���<���<���<���<���<���<���<���<���<���<ߐ�<Ր�<���<̐�<���<А�<���<А�<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<̐�<���<���<ɐ�<`   `   ���<���<�<o��<���<���<���<���<Ґ�<���<Ð�<���<���<���<���<o��<Ɛ�<���<���<���<ϐ�<���<ѐ�<���<`   `   
��<ϐ�<���<֐�<���<���<���<ϐ�<���<Ð�<Ԑ�<���<���<��<ѐ�<���<א�<��<ߐ�<���<ɐ�<Ő�<���<��<`   `   А�<Ӑ�<А�<��<���<���<Ґ�<���<���<���<ې�<���<���<��<��<Ӑ�<���<��<Ȑ�<��<Ґ�<��<���<��<`   `   ���<ߐ�<���<���<���<���<���<Ð�<���<���<���<ϐ�<���<���<ِ�<���<���<���<ݐ�<���<���<��<���<���<`   `   ���<���<���<���<���<���<Ð�<Ԑ�<ې�<���<���<���<���<���<���<���<
��<���<���<���<���<���<��<���<`   `   ���<���<���<���<���<���<���<���<���<ϐ�<���<���<���<���<���<Ր�<��<���<���<��<���<��<א�<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<А�<Ð�<��<Ð�<Ԑ�<���<���<���<`   `   ���<���<���<��<���<���<���<��<��<���<���<���<���<-��<��<���<��<��<��<���<���<��<.��<���<`   `   ���<ِ�<ː�<ѐ�<���<���<���<ѐ�<��<ِ�<���<���<���<��<���<ސ�<��<���<��<ސ�<���<��<���<���<`   `   ���<ސ�<���<b��<���<���<o��<���<Ӑ�<���<���<Ր�<���<���<ސ�<���<���<���<���<��<���<���<א�<���<`   `   ���<א�<Ȑ�<���<ߐ�<���<Ɛ�<א�<���<���<
��<��<А�<��<��<���<��<���<��<��<͐�<��<��<���<`   `   
��<���<���<��<Ր�<���<���<��<��<���<���<���<Ð�<��<���<���<���<���<��<�<���<���<���<���<`   `   Ԑ�<���<���<P��<���<���<���<ߐ�<Ȑ�<ݐ�<���<���<��<��<��<���<��<��<��<���<���<ݐ�<���<ߐ�<`   `   ���<ڐ�<���<~��<̐�<���<���<���<��<���<���<��<Ð�<���<ސ�<��<��<�<���<���<���<���<���<���<`   `   ���<ܐ�<���<ܐ�<���<̐�<ϐ�<ɐ�<Ґ�<���<���<���<Ԑ�<���<���<���<͐�<���<���<���<Đ�<ɐ�<ې�<̐�<`   `   ���<}��<���<���<А�<���<���<Ő�<��<��<���<��<���<��<��<���<��<���<ݐ�<���<ɐ�<���<���<ސ�<`   `   ���<���<���<͐�<���<���<ѐ�<���<���<���<��<א�<���<.��<���<א�<��<���<���<���<ې�<���<���<͐�<`   `   ֐�<ݐ�<��<ː�<А�<ɐ�<���<��<��<���<���<���<���<���<���<���<���<���<ߐ�<���<̐�<ސ�<͐�<ڐ�<`   `   ���<���<���<��<��<��<��<ݑ�<��<��<��<��<��<��<��<��<��<ݑ�<��<��<��<��< ��<���<`   `   ���<���<��<���<��<��<��<ϑ�<���<��<��<��<��<��<��<���<ӑ�<��<��<���<���<��<���<���<`   `   ���<��<0��<��<��<��<��<ґ�<Б�<��<��<��<��<��<̑�<ґ�<��<��<��<��<5��<��<���<��<`   `   ��<���<��<C��<��<���<%��<��<��<���<���<���<���<��<���<��<��<��<?��<���<���<��<��<��<`   `   ��<��<��<��<ő�<��<"��<	��<��<4��<��<4��<��<	��<,��<��<���<��<$��<��<��<��<��<��<`   `   ��<��<��<���<��<��<���<��<'��<��<��<-��<��<���<��<��<��<��<��<��<��<���<���< ��<`   `   ��<��<��<%��<"��<���<��<!��< ��<���<���<!��<$��<���<��<%��<��<��<��<���<��<ґ�<��<���<`   `   ݑ�<ϑ�<ґ�<��<	��<��<!��<"��<���< ��<%��<��<��<��<���<ˑ�<ӑ�<��<ܑ�<��<��<��<��<���<`   `   ��<���<Б�<��<��<'��< ��<���<:��<���<��<'��<��<��<ّ�<���<��<Ñ�<Ǒ�<��<��<��<�<Ñ�<`   `   ��<��<��<���<4��<��<���< ��<���<���<��<<��<���<ߑ�<��<��<��<ɑ�<��<ޑ�<���<��<ʑ�<��<`   `   ��<��<��<���<��<��<���<%��<��<��<��<���<��<��<��<��<��<���<!��<��<��<���<���<��<`   `   ��<��<��<���<4��<-��<!��<��<'��<<��<���<��<��<!��<��<Ց�<���<��<��<
��<��<��<֑�<��<`   `   ��<��<��<���<��<��<$��<��<��<���<��<��<��<���<Б�<���<��<���<���<���<��<���<̑�<���<`   `   ��<��<��<��<	��<���<���<��<��<ߑ�<��<!��<���<��<��<���<��<��<��<��<���<��<��<���<`   `   ��<��<̑�<���<,��<��<��<���<ّ�<��<��<��<Б�<��<֑�<Б�<��<��<���<Б�<ё�<��<ϑ�<��<`   `   ��<���<ґ�<��<��<��<%��<ˑ�<���<��<��<Ց�<���<���<Б�<��<��<ݑ�<��<ӑ�<���<���<֑�<ߑ�<`   `   ��<ӑ�<��<��<���<��<��<ӑ�<��<��<��<���<��<��<��<��<��<��<��<��<��<���<���<��<`   `   ݑ�<��<��<��<��<��<��<��<Ñ�<ɑ�<���<��<���<��<��<ݑ�<��<��<��<���<��<��<ʑ�<ɑ�<`   `   ��<��<��<?��<$��<��<��<ܑ�<Ǒ�<��<!��<��<���<��<���<��<��<��<���<��<"��<��<���<ܑ�<`   `   ��<���<��<���<��<��<���<��<��<ޑ�<��<
��<���<��<Б�<ӑ�<��<���<��<��<���<��<��<���<`   `   ��<���<5��<���<��<��<��<��<��<���<��<��<��<���<ё�<���<��<��<"��<���<���<��<��<��<`   `   ��<��<��<��<��<���<ґ�<��<��<��<���<��<���<��<��<���<���<��<��<��<��<ʑ�<���<��<`   `    ��<���<���<��<��<���<��<��<�<ʑ�<���<֑�<̑�<��<ϑ�<֑�<���<ʑ�<���<��<��<���<��<��<`   `   ���<���<��<��<��< ��<���<���<Ñ�<��<��<��<���<���<��<ߑ�<��<ɑ�<ܑ�<���<��<��<��<��<`   `   ���<\��<Q��<~��<^��<X��<F��<@��<a��<A��<%��<>��</��<>��<&��<A��<_��<@��<H��<X��<\��<~��<R��<\��<`   `   \��<P��<_��<5��<F��<@��<I��<f��<g��</��<��<%��<%��<��<.��<h��<f��<G��<?��<G��<5��<^��<Q��<]��<`   `   Q��<_��<���<-��<;��<'��<q��<p��<k��<f��<g��<S��<g��<f��<k��<p��<r��<'��<:��<-��<���<_��<P��<��<`   `   ~��<5��<-��<x��<��<F��<Y��<3��<[��<`��<.��<-��<`��<]��<3��<W��<G��<��<w��<,��<5��<��<3��<3��<`   `   ^��<F��<;��<��<-��<l��<��<,��<K��<"��<��<"��<J��<,��<��<l��<+��<��<=��<F��<]��<K��<J��<K��<`   `   X��<@��<'��<F��<l��<B��<F��<]��<6��<S��<S��<7��<]��<D��<B��<m��<G��<&��<?��<Y��<.��<Z��<Z��<.��<`   `   F��<I��<q��<Y��<��<F��<p��<��<B��<���<@��<��<r��<F��<��<Y��<r��<I��<F��<Z��<a��<i��<a��<Z��<`   `   @��<f��<p��<3��<,��<]��<��<���<W��<X��< ��<��<]��<-��<3��<o��<f��<A��<n��<��<:��<:��<��<o��<`   `   a��<g��<k��<[��<K��<6��<B��<W��<6��<W��<B��<6��<J��<[��<m��<g��<`��<���<w��<0��<!��<0��<w��<���<`   `   A��</��<f��<`��<"��<S��<���<X��<W��<���<S��<#��<`��<d��<.��<B��<���<���<J��<c��<c��<J��<���<���<`   `   %��<��<g��<.��<��<S��<@��< ��<B��<S��<��<.��<h��<��<$��<]��<C��<G��<S��<5��<R��<G��<C��<]��<`   `   >��<%��<S��<-��<"��<7��<��<��<6��<#��<.��<R��<%��<>��<���<j��<(��<~��<,��<-��<~��<(��<j��<���<`   `   /��<%��<g��<`��<J��<]��<r��<]��<J��<`��<h��<%��<.��<^��<x��<e��<l��<���<s��<���<m��<e��<x��<^��<`   `   >��<��<f��<]��<,��<D��<F��<-��<[��<d��<��<>��<^��<���<B��<k��<;��<���<���<:��<l��<C��<���<^��<`   `   &��<.��<k��<3��<��<B��<��<3��<m��<.��<$��<���<x��<B��<���<n��<I��<���<J��<n��<���<B��<x��<���<`   `   A��<h��<p��<W��<l��<m��<Y��<o��<g��<B��<]��<j��<e��<k��<n��<^��<f��<e��<]��<o��<l��<e��<j��<]��<`   `   _��<f��<r��<G��<+��<G��<r��<f��<`��<���<C��<(��<l��<;��<I��<f��<N��<f��<I��<;��<l��<(��<C��<���<`   `   @��<G��<'��<��<��<&��<I��<A��<���<���<G��<~��<���<���<���<e��<f��<���<���<���<~��<G��<���<���<`   `   H��<?��<:��<w��<=��<?��<F��<n��<w��<J��<S��<,��<s��<���<J��<]��<I��<���<t��<,��<T��<J��<v��<n��<`   `   X��<G��<-��<,��<F��<Y��<Z��<��<0��<c��<5��<-��<���<:��<n��<o��<;��<���<,��<4��<c��<1��<��<Y��<`   `   \��<5��<���<5��<]��<.��<a��<:��<!��<c��<R��<~��<m��<l��<���<l��<l��<~��<T��<c��< ��<:��<b��<.��<`   `   ~��<^��<_��<��<K��<Z��<i��<:��<0��<J��<G��<(��<e��<C��<B��<e��<(��<G��<J��<1��<:��<h��<Z��<M��<`   `   R��<Q��<P��<3��<J��<Z��<a��<��<w��<���<C��<j��<x��<���<x��<j��<C��<���<v��<��<b��<Z��<I��<3��<`   `   \��<]��<��<3��<K��<.��<Z��<o��<���<���<]��<���<^��<^��<���<]��<���<���<n��<Y��<.��<M��<3��<��<`   `   ���<���<���<���<���<���<���<Ô�<���<���<Ҕ�<���<ߔ�<���<Δ�<���<���<Ô�<���<���<���<���<���<���<`   `   ���<���<���<���<ʔ�<Ɣ�<ܔ�<���<���<Ɣ�<��<ה�<֔�<��<Ȕ�<���<���<��<Ȕ�<Ĕ�<���<���<��<���<`   `   ���<���<ה�<���<���<Ҕ�<x��<���<���<���<���<���<���<���<���<���<v��<Ҕ�<���<���<Ԕ�<���<���<Ӕ�<`   `   ���<���<���<���<ߔ�<ǔ�<p��<ϔ�<���<���<��<��<���<���<є�<v��<Ĕ�<ڔ�<���<��<���<���<۔�<ܔ�<`   `   ���<ʔ�<���<ߔ�<���<���<���<֔�<ǔ�<Ô�<��<Ô�<˔�<֔�<���<���<��<ߔ�<���<ʔ�<���<���<���<���<`   `   ���<Ɣ�<Ҕ�<ǔ�<���<Ҕ�<���<ɔ�<���<���<���<���<Ȕ�<���<Ԕ�<���<Ĕ�<֔�<Ȕ�<���<���<���<���<���<`   `   ���<ܔ�<x��<p��<���<���<���<ٔ�<�<���<Ȕ�<ٔ�<���<���<���<p��<w��<ܔ�<���<���<���<���<���<���<`   `   Ô�<���<���<ϔ�<֔�<ɔ�<ٔ�<��<���<���<��<ޔ�<Ȕ�<Д�<є�<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<ǔ�<���<�<���<O��<���<���<���<͔�<���<���<���<���<~��<���<���<��<���<���<~��<`   `   ���<Ɣ�<���<���<Ô�<���<���<���<���<���<���<���<���<���<Ȕ�<���<u��<���<���<��<��<���<���<x��<`   `   Ҕ�<��<���<��<��<���<Ȕ�<��<���<���<��<��<���<��<Ҕ�<���<���<���<���<���<���<���<���<���<`   `   ���<ה�<���<��<Ô�<���<ٔ�<ޔ�<���<���<��<���<֔�<���<o��<���<���<���<���<���<���<���<���<m��<`   `   ߔ�<֔�<���<���<˔�<Ȕ�<���<Ȕ�<͔�<���<���<֔�<��<���<�<���<���<Ɣ�<���<Ɣ�<���<���<Ĕ�<���<`   `   ���<��<���<���<֔�<���<���<Д�<���<���<��<���<���<��<���<|��<���<i��<k��<���<{��<���<��<���<`   `   Δ�<Ȕ�<���<є�<���<Ԕ�<���<є�<���<Ȕ�<Ҕ�<o��<�<���<���<���<���<���<���<���<���<���<�<o��<`   `   ���<���<���<v��<���<���<p��<���<���<���<���<���<���<|��<���<���<���<���<���<���<{��<���<���<���<`   `   ���<���<v��<Ĕ�<��<Ĕ�<w��<���<���<u��<���<���<���<���<���<���<v��<���<���<���<���<���<���<u��<`   `   Ô�<��<Ҕ�<ڔ�<ߔ�<֔�<ܔ�<���<~��<���<���<���<Ɣ�<i��<���<���<���<���<k��<Ɣ�<���<���<���<z��<`   `   ���<Ȕ�<���<���<���<Ȕ�<���<���<���<���<���<���<���<k��<���<���<���<k��<���<���<���<���<���<���<`   `   ���<Ĕ�<���<��<ʔ�<���<���<���<���<��<���<���<Ɣ�<���<���<���<���<Ɣ�<���<���<��<���<���<���<`   `   ���<���<Ԕ�<���<���<���<���<���<��<��<���<���<���<{��<���<{��<���<���<���<��<��<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<��<���<۔�<���<���<���<���<���<���<���<���<Ĕ�<��<�<���<���<���<���<���<���<���<���<۔�<`   `   ���<���<Ӕ�<ܔ�<���<���<���<���<~��<x��<���<m��<���<���<o��<���<u��<z��<���<���<���<���<۔�<ؔ�<`   `   ?��<4��<;��<���<&��<3��<��<L��<U��<\��<U��<��<=��<��<L��<\��<d��<L��<	��<3��<5��<���<2��<4��<`   `   4��<b��<:��<��<��<��<��<8��< ��<���<2��<��<��<7��<��<��<2��<��<��<���<��<D��<a��<.��<`   `   ;��<:��<$��<4��<��<=��<��<Y��<��<"��<)��<���<%��<"��<��<Y��<��<=��<��<4��<��<:��<B��<*��<`   `   ���<��<4��<��<��<E��<p��<G��<��<,��<��<��<+��<���<K��<|��<>��< ��<��<>��<��<���<��<��<`   `   &��<��<��<��<��<��<M��<��<-��<��<'��<��<7��<��<=��<��<���<��<��<��</��<(��<&��<(��<`   `   3��<��<=��<E��<��<L��<��<��<0��<��<��<'��<��<'��<P��<��<>��<G��<��<-��<p��<<��<;��<s��<`   `   ��<��<��<p��<M��<��<��<.��<���<��<��<.��<ܕ�<��<U��<p��<��<��<��<C��<&��<���<$��<C��<`   `   L��<8��<Y��<G��<��<��<.��<��</��<&��<��<9��<��<��<K��<c��<2��<F��<?��<M��<$��<'��<L��<9��<`   `   U��< ��<��<��<-��<0��<���</��<���</��<��<0��<:��<��<��< ��<a��<5��<g��<&��<��<&��<o��<5��<`   `   \��<���<"��<,��<��<��<��<&��</��<��<��<��<+��<,��<��<V��<!��<F��<A��<���<���<;��<E��<'��<`   `   U��<2��<)��<��<'��<��<��<��<��<��<7��<��<��<2��<V��<^��<=��<[��<&��<G��</��<[��<8��<^��<`   `   ��<��<���<��<��<'��<.��<9��<0��<��<��<��<��<��<���<;��<C��<��<Q��<K��<	��<J��<:��<���<`   `   =��<��<%��<+��<7��<��<ܕ�<��<:��<+��<��<��<C��<��<��<N��<'��< ��<:��< ��<$��<N��<$��<��<`   `   ��<7��<"��<���<��<'��<��<��<��<,��<2��<��<��<J��<6��<c��<���<5��<;��<���<_��<1��<I��<��<`   `   L��<��<��<K��<=��<P��<U��<K��<��<��<V��<���<��<6��<��<4��<e��<l��<Y��<4��<"��<6��<��<���<`   `   \��<��<Y��<|��<��<��<p��<c��< ��<V��<^��<;��<N��<c��<4��<��<D��<K��<��<0��<_��<O��<:��<b��<`   `   d��<2��<��<>��<���<>��<��<2��<a��<!��<=��<C��<'��<���<e��<D��<6��<D��<d��<���<*��<C��<:��<!��<`   `   L��<��<=��< ��<��<G��<��<F��<5��<F��<[��<��< ��<5��<l��<K��<D��<h��<;��<!��<	��<_��<E��<,��<`   `   	��<��<��<��<��<��<��<?��<g��<A��<&��<Q��<:��<;��<Y��<��<d��<;��<3��<Q��<%��<A��<q��<?��<`   `   3��<���<4��<>��<��<-��<C��<M��<&��<���<G��<K��< ��<���<4��<0��<���<!��<Q��<K��<���<��<L��<O��<`   `   5��<��<��<��</��<p��<&��<$��<��<���</��<	��<$��<_��<"��<_��<*��<	��<%��<���<��<$��<��<p��<`   `   ���<D��<:��<���<(��<<��<���<'��<&��<;��<[��<J��<N��<1��<6��<O��<C��<_��<A��<��<$��<	��<;��<��<`   `   2��<a��<B��<��<&��<;��<$��<L��<o��<E��<8��<:��<$��<I��<��<:��<:��<E��<q��<L��<��<;��<3��<��<`   `   4��<.��<*��<��<(��<s��<C��<9��<5��<'��<^��<���<��<��<���<b��<!��<,��<?��<O��<p��<��<��<4��<`   `   ���<���<���<��<�<���<֗�<���<���<���<���<���<���<���<���<���<Ɨ�<���<���<���<ؗ�<��<���<���<`   `   ���<���<���<ӗ�<���<ė�<���<���<���<}��<���<���<���<���<���<���<���<ŗ�<Η�<���<Η�<ŗ�<���<���<`   `   ���<���<X��<ɗ�<���<�<o��<���<��<��<ؗ�<���<ӗ�<��<��<���<h��<�< ��<ɗ�<O��<���<���<���<`   `   ��<ӗ�<ɗ�<֗�<���<՗�<���<j��<җ�<ߗ�<���<���<ޗ�<ŗ�<q��<×�<˗�<���<ߗ�<ؗ�<Η�<��<���<���<`   `   �<���<���<���<ϗ�<���<���<���<��<y��<���<y��<���<���<t��<���<��<���<ߗ�<���<З�<���<ȗ�<���<`   `   ���<ė�<�<՗�<���<���<ܗ�<��<���<���<���<���<��<��<���<���<˗�<ї�<Η�<���<���<���<���<���<`   `   ֗�<���<o��<���<���<ܗ�<ɗ�<ŗ�<���<��<���<ŗ�<���<ܗ�<���<���<j��<���<՗�<���<���<ϗ�<���<���<`   `   ���<���<���<j��<���<��<ŗ�<���<���<���<���<՗�<��<{��<q��<͗�<���<���<���<���<֗�<ۗ�<���<���<`   `   ���<���<��<җ�<��<���<���<���<՗�<���<���<���<���<җ�<˗�<���<�<���<���<���<՗�<���<���<���<`   `   ���<}��<��<ߗ�<y��<���<��<���<���<��<���<h��<ޗ�<��<���<z��<���<���<���<×�<���<���<���<���<`   `   ���<���<ؗ�<���<���<���<���<���<���<���<���<���<ʗ�<���<���<���<_��<���<���<���<���<���<V��<���<`   `   ���<���<���<���<y��<���<ŗ�<՗�<���<h��<���<��<���<���<��<���<���<���<���<���<���<���<���<��<`   `   ���<���<ӗ�<ޗ�<���<��<���<��<���<ޗ�<ʗ�<���<���<��<���<���<���<���<ʗ�<���<���<���<���<��<`   `   ���<���<��<ŗ�<���<��<ܗ�<{��<җ�<��<���<���<��<���<���<���<���<���<���<���<���<���<���<��<`   `   ���<���<��<q��<t��<���<���<q��<˗�<���<���<��<���<���<ė�<���<���<���<���<���<З�<���<���<��<`   `   ���<���<���<×�<���<���<���<͗�<���<z��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   Ɨ�<���<h��<˗�<��<˗�<j��<���<�<���<_��<���<���<���<���<���<���<���<���<���<���<���<Z��<���<`   `   ���<ŗ�<�<���<���<ї�<���<���<���<���<���<���<���<���<���<���<���<z��<���<���<���<���<���<���<`   `   ���<Η�< ��<ߗ�<ߗ�<Η�<՗�<���<���<���<���<���<ʗ�<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<ɗ�<ؗ�<���<���<���<���<���<×�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   ؗ�<Η�<O��<Η�<З�<���<���<֗�<՗�<���<���<���<���<���<З�<���<���<���<���<���<��<֗�<x��<���<`   `   ��<ŗ�<���<��<���<���<ϗ�<ۗ�<���<���<���<���<���<���<���<���<���<���<���<���<֗�<���<���<���<`   `   ���<���<���<���<ȗ�<���<���<���<���<���<V��<���<���<���<���<���<Z��<���<���<���<x��<���<ۗ�<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<��<��<��<��<���<���<���<���<���<���<���<���<���<`   `   ���<a��<4��<)��<Q��<4��<{��<+��<@��<K��<x��<]��<5��<]��<g��<K��<]��<+��<Z��<4��<n��<)��<#��<a��<`   `   a��<J��<h��<v��<��<��<���<x��<T��<��<q��<a��<_��<y��<���<D��<k��<���<+��<	��<o��<z��<I��<V��<`   `   4��<h��<"��<@��<=��<7��<$��<V��<]��<��<��<o��<ޘ�<��<c��<V��<��<7��<G��<@��<��<h��<?��<���<`   `   )��<v��<@��<&��<��<Q��<c��<A��<��<���<k��<r��<���<��<J��<x��<D��<���<3��<R��<o��<��<H��<I��<`   `   Q��<��<=��<��<r��<O��<���<��<h��<J��<���<J��<z��<��<f��<O��<���<��<��<��<c��<��<d��<��<`   `   4��<��<7��<Q��<O��<��<P��<(��<��<6��</��<���<&��<e��<��<9��<D��<I��<+��<*��<U��<[��<Z��<\��<`   `   {��<���<$��<c��<���<P��<ۘ�<[��<3��<��<J��<[��<Ș�<P��<���<c��<��<���<y��<���<V��<r��<P��<���<`   `   +��<x��<V��<A��<��<(��<[��<���<=��<.��<���<p��<&��<i��<J��<h��<k��< ��<L��<a��<7��<>��<_��<?��<`   `   @��<T��<]��<��<h��<��<3��<=��<r��<=��<%��<��<���<��<A��<T��<X��<Y��<k��<1��<4��<1��<x��<Y��<`   `   K��<��<��<���<J��<6��<��<.��<=��<(��</��<4��<���<1��<���<A��<���<���<?��<}��<v��<2��<��<���<`   `   x��<q��<��<k��<���</��<J��<���<%��</��<���<k��<Ә�<q��<y��<I��<_��<U��<H��<B��<\��<U��<S��<I��<`   `   ]��<a��<o��<r��<J��<���<[��<p��<��<4��<k��<���<_��<S��<7��<L��<���<���<��<��<���<���<K��<-��<`   `   5��<_��<ޘ�<���<z��<&��<Ș�<&��<���<���<Ә�<_��<A��<"��<K��<\��<X��<y��<���<y��<R��<\��<V��<"��<`   `   ]��<y��<��<��<��<e��<P��<i��<��<1��<q��<S��<"��<V��<��<I��<L��<c��<o��<Y��<B��<v��<U��<$��<`   `   g��<���<c��<J��<f��<��<���<J��<A��<���<y��<7��<K��<��<z��<]��<���<?��<m��<]��<���<��<K��<7��<`   `   K��<D��<V��<x��<O��<9��<c��<h��<T��<A��<I��<L��<\��<I��<]��<���<u��<���<���<T��<B��<^��<K��<P��<`   `   ]��<k��<��<D��<���<D��<��<k��<X��<���<_��<���<X��<L��<���<u��<��<u��<���<L��<]��<���<Y��<���<`   `   +��<���<7��<���<��<I��<���< ��<Y��<���<U��<���<y��<c��<?��<���<u��<5��<o��<{��<���<]��<��<I��<`   `   Z��<+��<G��<3��<��<+��<y��<L��<k��<?��<H��<��<���<o��<m��<���<���<o��<v��<��<H��<?��<{��<L��<`   `   4��<	��<@��<R��<��<*��<���<a��<1��<}��<B��<��<y��<Y��<]��<T��<L��<{��<��<I��<v��<"��<_��<���<`   `   n��<o��<��<o��<c��<U��<V��<7��<4��<v��<\��<���<R��<B��<���<B��<]��<���<H��<v��<K��<7��<B��<U��<`   `   )��<z��<h��<��<��<[��<r��<>��<1��<2��<U��<���<\��<v��<��<^��<���<]��<?��<"��<7��<���<Z��<��<`   `   #��<I��<?��<H��<d��<Z��<P��<_��<x��<��<S��<K��<V��<U��<K��<K��<Y��<��<{��<_��<B��<Z��<{��<H��<`   `   a��<V��<���<I��<��<\��<���<?��<Y��<���<I��<-��<"��<$��<7��<P��<���<I��<L��<���<U��<��<H��<���<`   `   ���<ۚ�<ܚ�<���<:��<��<Ӛ�<ۚ�<��<ʚ�<��<��<���<��<ޚ�<ʚ�<��<ۚ�<���<��<[��<���<ɚ�<ۚ�<`   `   ۚ�<0��<��<��< ��<К�<��<-��<њ�<��<��<��<��<!��<���<���<��<+��<ߚ�<��<���<,��<0��<К�<`   `   ܚ�<��<ʚ�<��<W��<%��<���<���<���<0��<��<���<ߚ�<0��<���<���<���<%��<`��<��<���<��<��<��<`   `   ���<��<��<
��<��<��<��<��<��<V��<���<��<R��<ޚ�<���<1��<���<��<��<(��<���<���<���<���<`   `   :��< ��<W��<��<��<Ě�<'��<֚�</��<$��<���<$��<D��<֚�<��<Ě�<:��<��<3��< ��<N��< ��<"��< ��<`   `   ��<К�<%��<��<Ě�<���<)��<��<��<��<��<��<��<@��<���<���<���<9��<ߚ�<ݚ�<#��<��<��<-��<`   `   Ӛ�<��<���<��<'��<)��<��<&��<���<.��<��<&��<��<)��<4��<��<���<��<Κ�<���<���<���<���<���<`   `   ۚ�<-��<���<��<֚�<��<&��<Ӛ�<��<ٚ�<˚�<=��<��<���<���<��<��<Ϛ�<��<���<��<��<���<ݚ�<`   `   ��<њ�<���<��</��<��<���<��<z��<��<��<��<K��<��<ؚ�<њ�<��<ך�<,��<��<��<��<<��<ך�<`   `   ʚ�<��<0��<V��<$��<��<.��<ٚ�<��<F��<��<��<R��<D��<���<���<��<Ț�<��<���<��<ܚ�<ǚ�<��<`   `   ��<��<��<���<���<��<��<˚�<��<��<֚�<���<Қ�<��<��<��<ݚ�<Κ�<��<��<��<Κ�<Κ�<��<`   `   ��<��<���<��<$��<��<&��<=��<��<��<���<��<��<��<��<��<��<ޚ�<��<���<՚�<���<��<ۚ�<`   `   ���<��<ߚ�<R��<D��<��<��<��<K��<R��<Қ�<��<��<��<��<��<���<՚�<��<՚�<���<��<#��<��<`   `   ��<!��<0��<ޚ�<֚�<@��<)��<���<��<D��<��<��<��<&��<њ�<��<*��<Ӛ�<��<:��<��<Ś�<%��<��<`   `   ޚ�<���<���<���<��<���<4��<���<ؚ�<���<��<��<��<њ�<њ�<ʚ�<��<��<��<ʚ�<��<њ�<��<��<`   `   ʚ�<���<���<1��<Ě�<���<��<��<њ�<���<��<��<��<��<ʚ�<���<��< ��<���<���<��<��<��<���<`   `   ��<��<���<���<:��<���<���<��<��<��<ݚ�<��<���<*��<��<��<���<��<���<*��<Ě�<��<ך�<��<`   `   ۚ�<+��<%��<��<��<9��<��<Ϛ�<ך�<Ț�<Κ�<ޚ�<՚�<Ӛ�<��< ��<��<ٚ�<��<ؚ�<՚�<֚�<ǚ�<ƚ�<`   `   ���<ߚ�<`��<��<3��<ߚ�<Κ�<��<,��<��<��<��<��<��<��<���<���<��<���<��<��<��<>��<��<`   `   ��<��<��<(��< ��<ݚ�<���<���<��<���<��<���<՚�<:��<ʚ�<���<*��<ؚ�<��<%��<��<���<���<��<`   `   [��<���<���<���<N��<#��<���<��<��<��<��<՚�<���<��<��<��<Ě�<՚�<��<��<���<��<���<#��<`   `   ���<,��<��<���< ��<��<���<��<��<ܚ�<Κ�<���<��<Ś�<њ�<��<��<֚�<��<���<��<��<��<��<`   `   ɚ�<0��<��<���<"��<��<���<���<<��<ǚ�<Κ�<��<#��<%��<��<��<ך�<ǚ�<>��<���<���<��<;��<���<`   `   ۚ�<К�<��<���< ��<-��<���<ݚ�<ך�<��<��<ۚ�<��<��<��<���<��<ƚ�<��<��<#��<��<���<-��<`   `   >��<�<���<Μ�<���<���<���<ڜ�<��<ל�<��<���<���<���<Ԝ�<ל�<��<ڜ�<Ӝ�<���<ڜ�<Μ�<���<�<`   `   �<���<Ɯ�<���<���<���<���<��<���<���<���<Ü�<���<���<���<���<Ϝ�<Ϝ�<���<q��<���<ڜ�<���<���<`   `   ���<Ɯ�<���<���<ݜ�<˜�<E��<ל�<��<М�<���<��<���<М�<��<ל�<@��<˜�<��<���<y��<Ɯ�<���<���<`   `   Μ�<���<���<F��<s��<ޜ�<Ϝ�<���<���<Ŝ�<���<Ŝ�<���<���<���<��<˜�<Z��<X��<͜�<���<Ü�<Ҝ�<ќ�<`   `   ���<���<ݜ�<s��<��<̜�<ќ�<n��<���<r��<|��<r��<���<n��<���<̜�<��<s��<���<���<̜�<���<���<���<`   `   ���<���<˜�<ޜ�<̜�<���<��<���<���<Ԝ�<͜�<���<���<���<���<���<˜�<ߜ�<���<���<���<���<���<���<`   `   ���<���<E��<Ϝ�<ќ�<��<���<ǜ�<���<
��<ʜ�<ǜ�<���<��<ܜ�<Ϝ�<D��<���<���<Ԝ�<���<)��<}��<Ԝ�<`   `   ڜ�<��<ל�<���<n��<���<ǜ�<f��<���<���<_��<ߜ�<���<U��<���<��<Ϝ�<Ϝ�<ٜ�<���<��<���<���<Ȝ�<`   `   ��<���<��<���<���<���<���<���<��<���<���<���<���<���<Ü�<���<���<���<Ӝ�<���<ɜ�<���<��<���<`   `   ל�<���<М�<Ŝ�<r��<Ԝ�<
��<���<���<"��<͜�<Y��<���<��<���<̜�<̜�<���<Ӝ�<���<���<���<���<ߜ�<`   `   ��<���<���<���<|��<͜�<ʜ�<_��<���<͜�<���<���<���<���<��<��<���<��<ʜ�<���<��<��<���<��<`   `   ���<Ü�<��<Ŝ�<r��<���<ǜ�<ߜ�<���<Y��<���<��<���<���<М�<̜�<��<��<М�<���<ڜ�<��<͜�<�<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<Ü�<���<Ŝ�<���<���<��<���<���<Ŝ�<ʜ�<Ü�<`   `   ���<���<М�<���<n��<���<��<U��<���<��<���<���<Ü�<���<���<��<��<���<���<��<��<���<���<Ȝ�<`   `   Ԝ�<���<��<���<���<���<ܜ�<���<Ü�<���<��<М�<���<���<��<ۜ�<���<՜�<Ϝ�<ۜ�<��<���<���<М�<`   `   ל�<���<ל�<��<̜�<���<Ϝ�<��<���<̜�<��<̜�<Ŝ�<��<ۜ�<���<��<��<���<͜�<��<ʜ�<͜�<��<`   `   ��<Ϝ�<@��<˜�<��<˜�<D��<Ϝ�<���<̜�<���<��<���<��<���<��<���<��<��<��<���<��<���<̜�<`   `   ڜ�<Ϝ�<˜�<Z��<s��<ߜ�<���<Ϝ�<���<���<��<��<���<���<՜�<��<��<ǜ�<���<���<ڜ�<��<���<���<`   `   Ӝ�<���<��<X��<���<���<���<ٜ�<Ӝ�<Ӝ�<ʜ�<М�<��<���<Ϝ�<���<��<���<���<М�<Ϝ�<Ӝ�<��<ٜ�<`   `   ���<q��<���<͜�<���<���<Ԝ�<���<���<���<���<���<���<��<ۜ�<͜�<��<���<М�<���<���<���<���<��<`   `   ڜ�<���<y��<���<̜�<���<���<��<ɜ�<���<��<ڜ�<���<��<��<��<���<ڜ�<Ϝ�<���<��<��<q��<���<`   `   Μ�<ڜ�<Ɯ�<Ü�<���<���<)��<���<���<���<��<��<Ŝ�<���<���<ʜ�<��<��<Ӝ�<���<��<A��<���<���<`   `   ���<���<���<Ҝ�<���<���<}��<���<��<���<���<͜�<ʜ�<���<���<͜�<���<���<��<���<q��<���<ǜ�<Ҝ�<`   `   �<���<���<ќ�<���<���<Ԝ�<Ȝ�<���<ߜ�<��<�<Ü�<Ȝ�<М�<��<̜�<���<ٜ�<��<���<���<Ҝ�<͜�<`   `   ���<m��<���<���<x��<���<���<M��<]��<{��<О�<���<���<���<���<{��<���<M��<n��<���<���<���<|��<m��<`   `   m��<l��<���<���<b��<a��<���<���<`��<t��<���<���<���<���<���<P��<���<���<u��<J��<���<���<n��<d��<`   `   ���<���<l��<֞�<Þ�<���<e��<���<���<���<K��<���<K��<���<���<���<c��<���<Ȟ�<֞�<e��<���<���<y��<`   `   ���<���<֞�<���<���<���<���<o��<���<o��<���<Ş�<i��<���<��<���<���<w��<���<��<���<���<���<���<`   `   x��<b��<Þ�<���<���<Y��<���<˞�<��<���<"��<���<���<˞�<x��<Y��<���<���<���<b��<���<c��<���<c��<`   `   ���<a��<���<���<Y��<e��<���<ʞ�<���<���<��<t��<Ğ�<���<t��<A��<���<Ξ�<u��<{��<���<���<���<���<`   `   ���<���<e��<���<���<���<��<���<}��<?��<���<���<ߝ�<���<���<���<g��<���<���<̞�<���<���<x��<̞�<`   `   M��<���<���<o��<˞�<ʞ�<���<��<���<���<��<Ğ�<Ğ�<���<��<˞�<���<D��<l��<���<L��<Y��<���<Y��<`   `   ]��<`��<���<���<��<���<}��<���<ƞ�<���<l��<���<��<���<z��<`��<{��<}��<���<s��<r��<s��<͞�<}��<`   `   {��<t��<���<o��<���<���<?��<���<���<V��<��<n��<i��<���<���<q��<���<���<e��<ޞ�<ў�<Q��<���<���<`   `   О�<���<K��<���<"��<��<���<��<l��<��<?��<���<>��<���<ʞ�<g��<Z��<���<N��<���<o��<���<C��<g��<`   `   ���<���<���<Ş�<���<t��<���<Ğ�<���<n��<���<���<���<���<i��<S��<���<���<S��<?��<���<���<U��<Y��<`   `   ���<���<K��<i��<���<Ğ�<ߝ�<Ğ�<��<i��<>��<���<���<|��<���<���<V��<���<��<���<N��<���<���<|��<`   `   ���<���<���<���<˞�<���<���<���<���<���<���<���<|��<���<���<r��<i��<t��<���<}��<e��<���<���<���<`   `   ���<���<���<��<x��<t��<���<��<z��<���<ʞ�<i��<���<���<x��<N��<���<m��<w��<N��<���<���<���<i��<`   `   {��<P��<���<���<Y��<A��<���<˞�<`��<q��<g��<S��<���<r��<N��<���<���<���<���<>��<e��<���<U��<l��<`   `   ���<���<c��<���<���<���<g��<���<{��<���<Z��<���<V��<i��<���<���<���<���<���<i��<\��<���<S��<���<`   `   M��<���<���<w��<���<Ξ�<���<D��<}��<���<���<���<���<t��<m��<���<���<]��<���<���<���<���<���<m��<`   `   n��<u��<Ȟ�<���<���<u��<���<l��<���<e��<N��<S��<��<���<w��<���<���<���<О�<S��<V��<e��<ɞ�<l��<`   `   ���<J��<֞�<��<b��<{��<̞�<���<s��<ޞ�<���<?��<���<}��<N��<>��<i��<���<S��<���<ў�<c��<���<��<`   `   ���<���<e��<���<���<���<���<L��<r��<ў�<o��<���<N��<e��<���<e��<\��<���<V��<ў�<���<L��<m��<���<`   `   ���<���<���<���<c��<���<���<Y��<s��<Q��<���<���<���<���<���<���<���<���<e��<c��<L��<���<���<K��<`   `   |��<n��<���<���<���<���<x��<���<͞�<���<C��<U��<���<���<���<U��<S��<���<ɞ�<���<m��<���<���<���<`   `   m��<d��<y��<���<c��<���<̞�<Y��<}��<���<g��<Y��<|��<���<i��<l��<���<m��<l��<��<���<K��<���<���<`   `   V��<t��<���<L��<���<|��<���<���<u��<q��<���<O��<|��<O��<k��<q��<���<���<Z��<|��<���<L��<t��<t��<`   `   t��<���<n��<���<y��<J��<���<���<g��<W��<u��<t��<l��<x��<g��<Y��<���<���<^��<d��<y��<��<���<m��<`   `   ���<n��<���<Q��<s��<a��<��<���<���<���<��<Z��<���<���<���<���<��<a��<t��<Q��<���<n��<���<���<`   `   L��<���<Q��<7��<q��<���<���<��<=��<���<<��<?��<���</��</��<���<q��<\��<K��<a��<y��<D��<g��<c��<`   `   ���<y��<s��<q��<_��<n��<���<(��<u��<)��<]��<)��<���<(��<p��<n��<���<q��<O��<y��<���<W��<Ǡ�<W��<`   `   |��<J��<a��<���<n��<���<���<���<D��<���<���<6��<���<���<���<Y��<q��<q��<^��<u��<l��<f��<i��<y��<`   `   ���<���<��<���<���<���<?��<f��<U��<���<f��<f��<3��<���<���<���<��<���<v��<P��<S��<P��<B��<P��<`   `   ���<���<���<��<(��<���<f��<l��<Y��<K��<h��<{��<���<��</��<���<���<���<0��<���<���<ɠ�<���<��<`   `   u��<g��<���<=��<u��<D��<U��<Y��<_��<Y��<D��<D��<���<=��<j��<g��<���<v��<���<|��<T��<|��<���<v��<`   `   q��<W��<���<���<)��<���<���<K��<Y��<à�<���<��<���<Ϡ�<g��<i��<���<���<6��<���<{��<!��<���<���<`   `   ���<u��<��<<��<]��<���<f��<h��<D��<���<u��<<��<v��<u��<v��<���<���<v��<���<��<���<v��<i��<���<`   `   O��<t��<Z��<?��<)��<6��<f��<{��<D��<��<<��<j��<l��<H��<|��<���<���<���<l��<X��<���<���<���<k��<`   `   |��<l��<���<���<���<���<3��<���<���<���<v��<l��<���<���<���<���<`��<���<l��<���<Y��<���<���<���<`   `   O��<x��<���</��<(��<���<���<��<=��<Ϡ�<u��<H��<���<A��<G��<���<���<V��<k��<Ӡ�<���<6��<E��<���<`   `   k��<g��<���</��<p��<���<���</��<j��<g��<v��<|��<���<G��<���<���<���<q��<���<���<Ơ�<G��<���<|��<`   `   q��<Y��<���<���<n��<Y��<���<���<g��<i��<���<���<���<���<���<e��<���<Ԡ�<y��<���<���<���<���<���<`   `   ���<���<��<q��<���<q��<��<���<���<���<���<���<`��<���<���<���<���<���<���<���<g��<���<{��<���<`   `   ���<���<a��<\��<q��<q��<���<���<v��<���<v��<���<���<V��<q��<Ԡ�<���<`��<k��<���<���<z��<���<h��<`   `   Z��<^��<t��<K��<O��<^��<v��<0��<���<6��<���<l��<l��<k��<���<y��<���<k��<P��<l��<���<6��<���<0��<`   `   |��<d��<Q��<a��<y��<u��<P��<���<|��<���<��<X��<���<Ӡ�<���<���<���<���<l��<��<{��<n��<���<d��<`   `   ���<y��<���<y��<���<l��<S��<���<T��<{��<���<���<Y��<���<Ơ�<���<g��<���<���<{��<o��<���<;��<l��<`   `   L��<��<n��<D��<W��<f��<P��<ɠ�<|��<!��<v��<���<���<6��<G��<���<���<z��<6��<n��<���<d��<i��<A��<`   `   t��<���<���<g��<Ǡ�<i��<B��<���<���<���<i��<���<���<E��<���<���<{��<���<���<���<;��<i��<٠�<g��<`   `   t��<m��<���<c��<W��<y��<P��<��<v��<���<���<k��<���<���<|��<���<���<h��<0��<d��<l��<A��<g��<���<`   `   ���<S��<L��<H��<_��<f��<���<���<;��<���<���<d��<}��<d��<���<���<Z��<���<���<f��<~��<H��<:��<S��<`   `   S��<1��<���<���<U��<8��<n��<Q��<k��<:��<:��<x��<p��<<��<K��<a��<<��<��<L��<D��<���<���<6��<N��<`   `   L��<���<f��<���<���<���<��<x��<���<<��<f��<���<m��<<��<���<x��<��<���<���<���<g��<���<L��<o��<`   `   H��<���<���<M��<c��<���<���<���<e��<���<���<���<���<[��<���<���<���<R��<a��<���<���<D��<L��<G��<`   `   _��<U��<���<c��<M��<H��<���<<��<��<t��<]��<t��<���<<��<j��<H��<s��<c��<s��<U��<r��<L��<���<L��<`   `   f��<8��<���<���<H��<��<X��<���<t��<���<���<i��<{��<h��</��<7��<���<���<L��<a��<��<d��<i��<���<`   `   ���<n��<��<���<���<X��<w��<���<V��<���<b��<���<o��<X��<���<���<��<n��<���<q��<T��<g��<A��<q��<`   `   ���<Q��<x��<���<<��<���<���<5��<n��<d��<3��<���<{��<+��<���<���<<��<���<Z��<T��<���<���<Y��<F��<`   `   ;��<k��<���<e��<��<t��<V��<n��<ˢ�<n��<G��<t��<���<e��<���<k��<U��<A��<���<K��<$��<K��<���<A��<`   `   ���<:��<<��<���<t��<���<���<d��<n��<���<���<b��<���<I��<K��<��<@��<`��<}��<L��<>��<i��<e��<U��<`   `   ���<:��<f��<���<]��<���<b��<3��<G��<���<o��<���<b��<:��<���<o��<B��<���<q��<A��<���<���<(��<o��<`   `   d��<x��<���<���<t��<i��<���<���<t��<b��<���<���<p��<_��<N��<T��<V��<y��<M��<9��<k��<k��<Y��<=��<`   `   }��<p��<m��<���<���<{��<o��<{��<���<���<b��<p��<���<���<s��<n��<��<p��<���<p��<��<n��<~��<���<`   `   d��<<��<<��<[��<<��<h��<X��<+��<e��<I��<:��<_��<���<V��<h��<���<y��<V��<j��<���<z��<W��<[��<���<`   `   ���<K��<���<���<j��</��<���<���<���<K��<���<N��<s��<h��<���<G��<x��<s��<O��<G��<���<h��<e��<N��<`   `   ���<a��<x��<���<H��<7��<���<���<k��<��<o��<T��<n��<���<G��<��<[��<p��<���<7��<z��<w��<Y��<p��<`   `   Z��<<��<��<���<s��<���<��<<��<U��<@��<B��<V��<��<y��<x��<[��<��<[��<u��<y��<��<V��<<��<@��<`   `   ���<��<���<R��<c��<���<n��<���<A��<`��<���<y��<p��<V��<s��<p��<[��<b��<j��<x��<k��<���<e��<7��<`   `   ���<L��<���<a��<s��<L��<���<Z��<���<}��<q��<M��<���<j��<O��<���<u��<j��<y��<M��<~��<}��<���<Z��<`   `   f��<D��<���<���<U��<a��<q��<T��<K��<L��<A��<9��<p��<���<G��<7��<y��<x��<M��<B��<>��<A��<Y��<���<`   `   ~��<���<g��<���<r��<��<T��<���<$��<>��<���<k��<��<z��<���<z��<��<k��<~��<>��<=��<���<>��<��<`   `   H��<���<���<D��<L��<d��<g��<���<K��<i��<���<k��<n��<W��<h��<w��<V��<���<}��<A��<���<w��<i��<;��<`   `   :��<6��<L��<L��<���<i��<A��<Y��<���<e��<(��<Y��<~��<[��<e��<Y��<<��<e��<���<Y��<>��<i��<���<L��<`   `   S��<N��<o��<G��<L��<���<q��<F��<A��<U��<o��<=��<���<���<N��<p��<@��<7��<Z��<���<��<;��<L��<|��<`   `   ���<d��<���<���<R��<Z��<c��<X��<e��<q��<���<���<:��<���<���<q��<~��<X��<E��<Z��<k��<���<z��<d��<`   `   d��<6��<z��<V��<E��<4��<s��<���<z��<W��<Ĥ�<��<v��<ä�<f��<s��<���<��<F��<9��<I��<���<<��<a��<`   `   ���<z��<���<v��<���<���<f��<\��<��<V��<D��<S��<M��<V��<v��<\��<m��<���<���<v��<��<z��<���<���<`   `   ���<V��<v��<K��<,��<���<:��<A��<w��<X��<a��<`��<O��<q��<P��<E��<���< ��<]��<��<I��<���<���<z��<`   `   R��<E��<���<,��<T��<Z��<���<���<v��<s��<���<s��<���<���<m��<Z��<s��<,��<���<E��<a��<a��<\��<a��<`   `   Z��<4��<���<���<Z��<q��<���<T��<c��<A��<B��<]��<K��<���<���<N��<���<���<F��<X��<���<_��<e��<���<`   `   c��<s��<f��<:��<���<���<��<���<i��<'��<o��<���<��<���<���<:��<p��<s��<S��<���<t��<���<a��<���<`   `   X��<���<\��<A��<���<T��<���<���<\��<V��<���<���<K��<���<P��<e��<���<V��<u��<G��<Y��<f��<M��<c��<`   `   e��<z��<��<w��<v��<c��<i��<\��<|��<\��<]��<c��<���<w��<f��<z��<z��<���<���<s��<���<s��<���<���<`   `   q��<W��<V��<X��<s��<A��<'��<V��<\��<2��<B��<g��<O��<_��<f��<o��<���<}��<z��<���<��<h��<���<���<`   `   ���<Ĥ�<D��<a��<���<B��<o��<���<]��<B��<���<a��<D��<Ĥ�<���<{��<���<c��<Y��<d��<y��<c��<t��<{��<`   `   ���<��<S��<`��<s��<]��<���<���<c��<g��<a��<\��<v��<���<?��<v��<���<���<���<w��<���<Ƥ�<|��<0��<`   `   :��<v��<M��<O��<���<K��<��<K��<���<O��<D��<v��<E��<t��<���<Ĥ�<i��<���<��<���<d��<Ĥ�<���<t��<`   `   ���<ä�<V��<q��<���<���<���<���<w��<_��<Ĥ�<���<t��<���<���<���<���<D��<V��<���<���<{��<���<}��<`   `   ���<f��<v��<P��<m��<���<���<P��<f��<f��<���<?��<���<���<K��<���<ۤ�<���<���<���<h��<���<{��<?��<`   `   q��<s��<\��<E��<Z��<N��<:��<e��<z��<o��<{��<v��<Ĥ�<���<���<Τ�<¤�<դ�<��<u��<���<ͤ�<|��<{��<`   `   ~��<���<m��<���<s��<���<p��<���<z��<���<���<���<i��<���<ۤ�<¤�<#��<¤�<٤�<���<n��<���<���<���<`   `   X��<��<���< ��<,��<���<s��<V��<���<}��<c��<���<���<D��<���<դ�<¤�<s��<V��<���<���<b��<���<��<`   `   E��<F��<���<]��<���<F��<S��<u��<���<z��<Y��<���<��<V��<���<��<٤�<V��<Ҥ�<���<g��<z��<���<u��<`   `   Z��<9��<v��<��<E��<X��<���<G��<s��<���<d��<w��<���<���<���<u��<���<���<���<c��<��<l��<M��<���<`   `   k��<I��<��<I��<a��<���<t��<Y��<���<��<y��<���<d��<���<h��<���<n��<���<g��<��<���<Y��<c��<���<`   `   ���<���<z��<���<a��<_��<���<f��<s��<h��<c��<Ƥ�<Ĥ�<{��<���<ͤ�<���<b��<z��<l��<Y��<���<e��<T��<`   `   z��<<��<���<���<\��<e��<a��<M��<���<���<t��<|��<���<���<{��<|��<���<���<���<M��<c��<e��<c��<���<`   `   d��<a��<���<z��<a��<���<���<c��<���<���<{��<0��<t��<}��<?��<{��<���<��<u��<���<���<T��<���<���<`   `   \��<���<s��<{��<���<���<���<a��<r��<R��<e��<���<a��<���<[��<R��<���<a��<���<���<���<{��<i��<���<`   `   ���<���<���<���<���<���<���<��<���<X��<���<���<���<���<e��<���<զ�<���<���<���<���<���<���<���<`   `   s��<���<d��<���<���<A��<o��<���<���<٦�<���<���<���<٦�<���<���<x��<A��<���<���<k��<���<m��<d��<`   `   {��<���<���<���<n��<���<���<Q��<���<���<���<���<���<���<]��<���<���<h��<���<���<���<|��<]��<W��<`   `   ���<���<���<n��<���<���<���<���<s��<���<���<���<~��<���<���<���<Ц�<n��<���<���<���<���<���<���<`   `   ���<���<A��<���<���<o��<���<���<���<���<���<���<���<���<{��<���<���<E��<���<���<`��<s��<y��<l��<`   `   ���<���<o��<���<���<���<x��<���<���<צ�<���<���<z��<���<���<���<z��<���<���<���<z��<���<i��<���<`   `   a��<��<���<Q��<���<���<���<r��<���<���<u��<���<���<���<]��<���<զ�<a��<���<���<���<���<���<���<`   `   r��<���<���<���<s��<���<���<���<��<���<���<���<���<���<���<���<���<���<���<h��<C��<h��<���<���<`   `   R��<X��<٦�<���<���<���<צ�<���<���<ަ�<���<���<���<ަ�<e��<R��<���<j��<W��<|��<q��<I��<q��<̦�<`   `   e��<���<���<���<���<���<���<u��<���<���<���<���<���<���<X��<���<���<z��<���<t��<���<z��<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<Ħ�<���<z��<���<���<���<���<`   `   a��<���<���<���<~��<���<z��<���<���<���<���<���<h��<���<���<q��<a��<���<���<���<]��<q��<���<���<`   `   ���<���<٦�<���<���<���<���<���<���<ަ�<���<���<���<���<d��<���<���<l��<{��<Ŧ�<���<W��<���<Ȧ�<`   `   [��<e��<���<]��<���<{��<���<]��<���<e��<X��<���<���<d��<���<���<���<s��<���<���<¦�<d��<���<���<`   `   R��<���<���<���<���<���<���<���<���<R��<���<���<q��<���<���<6��<���<���<E��<���<���<y��<���<���<`   `   ���<զ�<x��<���<Ц�<���<z��<զ�<���<���<���<���<a��<���<���<���<r��<���<���<���<d��<���<���<���<`   `   a��<���<A��<h��<n��<E��<���<a��<���<j��<z��<Ħ�<���<l��<s��<���<���<f��<{��<���<���<w��<q��<���<`   `   ���<���<���<���<���<���<���<���<���<W��<���<���<���<{��<���<E��<���<{��<���<���<���<W��<���<���<`   `   ���<���<���<���<���<���<���<���<h��<|��<t��<z��<���<Ŧ�<���<���<���<���<���<r��<q��<f��<���<���<`   `   ���<���<k��<���<���<`��<z��<���<C��<q��<���<���<]��<���<¦�<���<d��<���<���<q��<Q��<���<n��<`��<`   `   {��<���<���<|��<���<s��<���<���<h��<I��<z��<���<q��<W��<d��<y��<���<w��<W��<f��<���<Ȧ�<y��<���<`   `   i��<���<m��<]��<���<y��<i��<���<���<q��<���<���<���<���<���<���<���<q��<���<���<n��<y��<���<]��<`   `   ���<���<d��<W��<���<l��<���<���<���<̦�<���<���<���<Ȧ�<���<���<���<���<���<���<`��<���<]��<h��<`   `   P��<ʨ�<���<���<���<���<��<���<���<���<��<ʨ�<ʨ�<ʨ�<��<���<���<���<ݨ�<���<���<���<���<ʨ�<`   `   ʨ�<���<���<˨�<{��<���<֨�<���<���<ڨ�<���<��<ި�<���<��<���<���<֨�<���<z��<è�<���<���<ͨ�<`   `   ���<���<ܨ�<���<���<���<���<���<���<���<}��<٨�<���<���<���<���<���<���<���<���<��<���<���<��<`   `   ���<˨�<���<���<��<���<��<���<���<Ũ�<���<���<���<���<Ȩ�<��<���< ��<���<���<è�<���<���<���<`   `   ���<{��<���<��<���<���<���<���<���<���<���<���<¨�<���<��<���<���<��<���<{��<���<ݨ�<��<ݨ�<`   `   ���<���<���<���<���<C��<���<��<���<r��<v��<���<ڨ�<���<L��<���<���<���<���<���<���<���<���<ƨ�<`   `   ��<֨�<���<��<���<���<ݨ�<ɨ�<���<���<���<ɨ�<��<���<��<��<���<֨�<ܨ�<���<���<���<���<���<`   `   ���<���<���<���<���<��<ɨ�<j��<���<���<n��<ʨ�<ڨ�<���<Ȩ�<���<���<���<���<���<Ш�<ب�<���<���<`   `   ���<���<���<���<���<���<���<���<Ҩ�<���<���<���<Ĩ�<���<���<���<���<���<��<��<���<��<��<���<`   `   ���<ڨ�<���<Ũ�<���<r��<���<���<���<���<v��<���<���<���<��<���<̨�<���<���<��<��<��<���<֨�<`   `   ��<���<}��<���<���<v��<���<n��<���<v��<���<���<���<���<��<Ψ�<���<���<��<ب�<��<���<���<Ψ�<`   `   ʨ�<��<٨�<���<���<���<ɨ�<ʨ�<���<���<���<٨�<ި�<ͨ�<��<���<٨�<��<���<���<��<��<���<��<`   `   ʨ�<ި�<���<���<¨�<ڨ�<��<ڨ�<Ĩ�<���<���<ި�<Ψ�<Ǩ�<��<ܨ�<���<���<���<���<���<ܨ�<��<Ǩ�<`   `   ʨ�<���<���<���<���<���<���<���<���<���<���<ͨ�<Ǩ�<���<���<���<��<��<��<���<���<��<���<ͨ�<`   `   ��<��<���<Ȩ�<��<L��<��<Ȩ�<���<��<��<��<��<���<���<���<��< ��<��<���<
��<���<٨�<��<`   `   ���<���<���<��<���<���<��<���<���<���<Ψ�<���<ܨ�<���<���<���<��<��<���<���<���<��<���<ʨ�<`   `   ���<���<���<���<���<���<���<���<���<̨�<���<٨�<���<��<��<��< ��<��<��<��<���<٨�<���<̨�<`   `   ���<֨�<���< ��<��<���<֨�<���<���<���<���<��<���<��< ��<��<��<���<��<Ũ�<��<��<���<���<`   `   ݨ�<���<���<���<���<���<ܨ�<���<��<���<��<���<���<��<��<���<��<��<��<���<��<���<ߨ�<���<`   `   ���<z��<���<���<{��<���<���<���<��<��<ب�<���<���<���<���<���<��<Ũ�<���<ը�<��<��<���<���<`   `   ���<è�<��<è�<���<���<���<Ш�<���<��<��<��<���<���<
��<���<���<��<��<��<���<Ш�<���<���<`   `   ���<���<���<���<ݨ�<���<���<ب�<��<��<���<��<ܨ�<��<���<��<٨�<��<���<��<Ш�<���<���<ܨ�<`   `   ���<���<���<���<��<���<���<���<��<���<���<���<��<���<٨�<���<���<���<ߨ�<���<���<���<��<���<`   `   ʨ�<ͨ�<��<���<ݨ�<ƨ�<���<���<���<֨�<Ψ�<��<Ǩ�<ͨ�<��<ʨ�<̨�<���<���<���<���<ܨ�<���<��<`   `   ���<ݪ�<���<��<��<ڪ�<��<��<��<��<	��<��<��<��<	��<��<��<��<��<ڪ�<��<��<���<ݪ�<`   `   ݪ�<ߪ�<˪�<��<��<��<���<��<���<��<��<��<��<��<��< ��<
��<���<��<��<��<Ǫ�<��<��<`   `   ���<˪�<��<��<��<��<��<��<���<��<���<��<���<��<��<��<	��<��<��<��<��<˪�<���<ݪ�<`   `   ��<��<��<���<٪�<��<��<ɪ�<��<#��<���<���<��<
��<ͪ�<��<��<ݪ�<���<��<��<��<۪�<ת�<`   `   ��<��<��<٪�<���<��<��<��<��<��<)��<��<��<��<��<��<���<٪�<��<��<��<ت�<���<ت�<`   `   ڪ�<��<��<��<��<Q��<��<ת�<��<��<��<��<Ӫ�<��<U��<��<��<��<��<ު�<5��<֪�<ڪ�<9��<`   `   ��<���<��<��<��<��<ʪ�<��<&��<��<��<��<Ҫ�<��<��<��<	��<���<��<��</��<��<'��<��<`   `   ��<��<��<ɪ�<��<ת�<��<;��<��<��<?��<��<Ӫ�<��<ͪ�<��<
��< ��<��<̪�<��<��<Ъ�<��<`   `   ��<���<���<��<��<��<&��<��<���<��<&��<��<��<��<���<���<��<$��<��<���<��<���<��<$��<`   `   ��<��<��<#��<��<��<��<��<��<��<��<��<��<
��<��<���<��<��<Ϊ�< ��<���<ʪ�<��<��<`   `   	��<��<���<���<)��<��<��<?��<&��<��<!��<���<���<��<��<ɪ�<(��<��<���<���<���<��< ��<ɪ�<`   `   ��<��<��<���<��<��<��<��<��<��<���<��<��<��<��<��<J��<��<��<��<��<N��<	��<ު�<`   `   ��<��<���<��<��<Ӫ�<Ҫ�<Ӫ�<��<��<���<��<��<��<��<-��<#��<!��<5��<!��<#��<-��<��<��<`   `   ��<��<��<
��<��<��<��<��<��<
��<��<��<��<��<���<���<��<Ǫ�<̪�<��<��<���<��<��<`   `   	��<��<��<ͪ�<��<U��<��<ͪ�<���<��<��<��<��<���<ʪ�<��<��<���<��<��<Ҫ�<���<
��<��<`   `   ��< ��<��<��<��<��<��<��<���<���<ɪ�<��<-��<���<��<���<���<��<���<��<��<1��<	��<Ū�<`   `   ��<
��<	��<��<���<��<	��<
��<��<��<(��<J��<#��<��<��<���<���<���<��<��<#��<J��<(��<��<`   `   ��<���<��<ݪ�<٪�<��<���< ��<$��<��<��<��<!��<Ǫ�<���<��<���<���<̪�<%��<��<ު�<��<(��<`   `   ��<��<��<���<��<��<��<��<��<Ϊ�<���<��<5��<̪�<��<���<��<̪�<-��<��<���<Ϊ�<ު�<��<`   `   ڪ�<��<��<��<��<ު�<��<̪�<���< ��<���<��<!��<��<��<��<��<%��<��<���<���<���<Ъ�<��<`   `   ��<��<��<��<��<5��</��<��<��<���<���<��<#��<��<Ҫ�<��<#��<��<���<���<��<��</��<5��<`   `   ��<Ǫ�<˪�<��<ت�<֪�<��<��<���<ʪ�<��<N��<-��<���<���<1��<J��<ު�<Ϊ�<���<��<��<ڪ�<ܪ�<`   `   ���<��<���<۪�<���<ڪ�<'��<Ъ�<��<��< ��<	��<��<��<
��<	��<(��<��<ު�<Ъ�</��<ڪ�<���<۪�<`   `   ݪ�<��<ݪ�<ת�<ت�<9��<��<��<$��<��<ɪ�<ު�<��<��<��<Ū�<��<(��<��<��<5��<ܪ�<۪�<٪�<`   `   ���<'��<B��<L��<���<P��<@��<@��<*��<E��<\��<n��<G��<n��<b��<E��< ��<@��<K��<P��<��<L��<G��<'��<`   `   '��<K��</��<��<f��<-��<���<P��<X��<��<W��<<��<;��<S��<��<^��<S��<���<*��<o��<��<(��<M��<,��<`   `   B��</��<��<O��<Q��<.��<]��<���<a��<3��<z��<J��<~��<3��<\��<���<c��<.��<K��<O��<��</��<;��<¬�<`   `   L��<��<O��<6��<<��<U��<���<[��<j��<3��<A��<=��<3��<q��<Z��<���<X��<D��<4��<H��<��<Q��<a��<_��<`   `   ���<f��<Q��<<��<���<S��<ެ�<w��<.��<��<<��<��<(��<w��<��<S��<���<<��<[��<f��<���<)��<y��<)��<`   `   P��<-��<.��<U��<S��<��<A��<s��<E��<E��<I��<L��<r��<8��<��<\��<X��<'��<*��<U��<��<X��<Y��<��<`   `   @��<���<]��<���<ެ�<A��<X��<1��<<��<���<1��<1��<a��<A��<׬�<���<b��<���<>��<=��<.��<Z��<-��<=��<`   `   @��<P��<���<[��<w��<s��<1��<3��<,��<2��<7��<(��<r��<���<Z��<���<S��<E��<f��<K��<L��<L��<M��<i��<`   `   *��<X��<a��<j��<.��<E��<<��<,��<L��<,��<@��<E��<&��<j��<j��<X��<"��<9��<k��<���<F��<���<f��<9��<`   `   E��<��<3��<3��<��<E��<���<2��<,��<���<I��<��<3��<+��<��<J��<Q��<]��<���<l��<m��<���<_��<N��<`   `   \��<W��<z��<A��<<��<I��<1��<7��<@��<I��<0��<A��<���<W��<Y��<��<���<p��<���<���<���<p��<���<��<`   `   n��<<��<J��<=��<��<L��<1��<(��<E��<��<A��<C��<;��<s��<���<`��<A��<p��<���<���<q��<>��<b��<���<`   `   G��<;��<~��<3��<(��<r��<a��<r��<&��<3��<���<;��<C��<���<y��<2��<x��<���<Y��<���<z��<2��<v��<���<`   `   n��<S��<3��<q��<w��<8��<A��<���<j��<+��<W��<s��<���<���<|��<���<���<���<���<���<���<~��<���<���<`   `   b��<��<\��<Z��<��<��<׬�<Z��<j��<��<Y��<���<y��<|��<ԭ�<}��<}��<���<���<}��<ҭ�<|��<w��<���<`   `   E��<^��<���<���<S��<\��<���<���<X��<J��<��<`��<2��<���<}��<F��<���<���<C��<~��<���<3��<b��<{��<`   `    ��<S��<c��<X��<���<X��<b��<S��<"��<Q��<���<A��<x��<���<}��<���<���<���<~��<���<v��<A��<���<Q��<`   `   @��<���<.��<D��<<��<'��<���<E��<9��<]��<p��<p��<���<���<���<���<���<���<���<���<q��<l��<_��<@��<`   `   K��<*��<K��<4��<[��<*��<>��<f��<k��<���<���<���<Y��<���<���<C��<~��<���<[��<���<���<���<b��<f��<`   `   P��<o��<O��<H��<f��<U��<=��<K��<���<l��<���<���<���<���<}��<~��<���<���<���<���<m��<���<M��<5��<`   `   ��<��<��<��<���<��<.��<L��<F��<m��<���<q��<z��<���<ҭ�<���<v��<q��<���<m��<>��<L��<4��<��<`   `   L��<(��</��<Q��<)��<X��<Z��<L��<���<���<p��<>��<2��<~��<|��<3��<A��<l��<���<���<L��<Q��<Y��<1��<`   `   G��<M��<;��<a��<y��<Y��<-��<M��<f��<_��<���<b��<v��<���<w��<b��<���<_��<b��<M��<4��<Y��<o��<a��<`   `   '��<,��<¬�<_��<)��<��<=��<i��<9��<N��<��<���<���<���<���<{��<Q��<@��<f��<5��<��<1��<a��<���<`   `   ���<|��<���<���<���<��<���<��<ۯ�<��<���<���<��<���<ů�<��<ɯ�<��<ԯ�<��<���<���<���<|��<`   `   |��<d��<���<z��<v��<���<���<y��<���<��<Ư�<���<���<ï�<گ�<���<���<���<���<���<���<���<d��<���<`   `   ���<���<ԯ�<}��<]��<���<˯�<���<~��<���<��<���<��<���<}��<���<ͯ�<���<Z��<}��<د�<���<���<���<`   `   ���<z��<}��<���<���<���<���<��<���<���<ͯ�<ʯ�<���<���<ۯ�<���<���<���<���<s��<���<���<���<���<`   `   ���<v��<]��<���<`��<���<į�<���<���<̯�<���<̯�<|��<���<ׯ�<���<J��<���<q��<v��<���<���<t��<���<`   `   ��<���<���<���<���<ί�<���<���<կ�<���<���<ݯ�<���<��<ǯ�<˯�<���<���<���<��<���<���<���<���<`   `   ���<���<˯�<���<į�<���<���<���<���<���<���<���<���<���<���<���<˯�<���<ï�<���<���<���<���<���<`   `   ��<y��<���<��<���<���<���<���<̯�<կ�<���<���<���<���<ۯ�<y��<���<��<���<���<Ư�<���<���<���<`   `   ۯ�<���<~��<���<���<կ�<���<̯�<��<̯�<ǯ�<կ�<x��<���<���<���<̯�<���<���<į�<���<į�<���<���<`   `   ��<��<���<���<̯�<���<���<կ�<̯�<���<���<ٯ�<���<���<گ�<��<���<���<���<s��<y��<¯�<���<���<`   `   ���<Ư�<��<ͯ�<���<���<���<���<ǯ�<���<���<ͯ�<��<Ư�<���<���<���<ѯ�<��<���<د�<ѯ�<ï�<���<`   `   ���<���<���<ʯ�<̯�<ݯ�<���<���<կ�<ٯ�<ͯ�<���<���<���<���<��<¯�<߯�<���<���<��<���<��<���<`   `   ��<���<��<���<|��<���<���<���<x��<���<��<���<د�<���<ܯ�< ��<��<ܯ�<���<ܯ�<��< ��<կ�<���<`   `   ���<ï�<���<���<���<��<���<���<���<���<Ư�<���<���<���<ï�<ۯ�<į�<���<��<���<��<˯�<���<���<`   `   ů�<گ�<}��<ۯ�<ׯ�<ǯ�<���<ۯ�<���<گ�<���<���<ܯ�<ï�<��<��<���<��<���<��<��<ï�<��<���<`   `   ��<���<���<���<���<˯�<���<y��<���<��<���<��< ��<ۯ�<��<߯�<ί�<į�<֯�<���<��<���<��<���<`   `   ɯ�<���<ͯ�<���<J��<���<˯�<���<̯�<���<���<¯�<��<į�<���<ί�<��<ί�<���<į�<���<¯�<���<���<`   `   ��<���<���<���<���<���<���<��<���<���<ѯ�<߯�<ܯ�<���<��<į�<ί�<���<��<گ�<��<ί�<���<���<`   `   ԯ�<���<Z��<���<q��<���<ï�<���<���<���<��<���<���<��<���<֯�<���<��<���<���<��<���<���<���<`   `   ��<���<}��<s��<v��<��<���<���<į�<s��<���<���<ܯ�<���<��<���<į�<گ�<���<���<y��<ͯ�<���<x��<`   `   ���<���<د�<���<���<���<���<Ư�<���<y��<د�<��<��<��<��<��<���<��<��<y��<���<Ư�<���<���<`   `   ���<���<���<���<���<���<���<���<į�<¯�<ѯ�<���< ��<˯�<ï�<���<¯�<ί�<���<ͯ�<Ư�<���<���<���<`   `   ���<d��<���<���<t��<���<���<���<���<���<ï�<��<կ�<���<��<��<���<���<���<���<���<���<h��<���<`   `   |��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<x��<���<���<���<���<`   `   |��<���<���<��<#��<��<���<��<,��<	��<��<X��<���<X��<��<	��<��<��<ұ�<��<��<��<��<���<`   `   ���<ձ�<ϱ�<���<��<��<��<��<,��<f��<��<=��<C��<��<Y��<5��<��<��<
��<��<��<ñ�<ұ�<��<`   `   ���<ϱ�<F��<���<��<#��<L��<���<-��<7��<$��<��< ��<7��<1��<���<J��<#��<��<���<G��<ϱ�<���<E��<`   `   ��<���<���<N��<=��<��<	��<.��<5��<F��<��<��<L��<?��<!��<���<��<L��<>��<��<��<��<߱�<��<`   `   #��<��<��<=��<��<��<��< ��<��<6��<��<6��<��< ��<��<��<ı�<=��<��<��<��<��<ı�<��<`   `   ��<��<#��<��<��<;��<��<���<��<���<���<��< ��<���<.��<$��<��<��<
��<���<��<��<��<��<`   `   ���<��<L��<	��<��<��<Y��<��<#��<��<��<��<b��<��< ��<	��<G��<��<���<��<G��<��<V��<��<`   `   ��<��<���<.��< ��<���<��<��<���<��<��<���< ��<��<!��<��<��<#��<��<Q��<��<��<N��<"��<`   `   ,��<,��<-��<5��<��<��<#��<���<Z��<���</��<��<���<5��<G��<,��<��<^��<��<?��<|��<?��<��<^��<`   `   	��<f��<7��<F��<6��<���<��<��<���<��<���<F��<L��<*��<Y��<��<!��<���<<��<{��<���<L��<���<��<`   `   ��<��<$��<��<��<���<��<��</��<���<ڱ�<��<*��<��<��<��<o��<^��<S��<���<8��<^��<���<��<`   `   X��<=��<��<��<6��<��<��<���<��<F��<��<��<C��<]��<Z��<h��<A��<:��<���<���<E��<0��<e��<g��<`   `   ���<C��< ��<L��<��< ��<b��< ��<���<L��<*��<C��<���<c��<���<}��<���<���<���<���<���<}��<���<c��<`   `   X��<��<7��<?��< ��<���<��<��<5��<*��<��<]��<c��<���<���<4��<f��<���<���<V��<?��<���<���<]��<`   `   ��<Y��<1��<!��<��<.��< ��<!��<G��<Y��<��<Z��<���<���<-��<���<���<X��<���<���<��<���<���<Z��<`   `   	��<5��<���<���<��<$��<	��<��<,��<��<��<h��<}��<4��<���<@��<���<���<0��<Ų�<?��<v��<e��<	��<`   `   ��<��<J��<��<ı�<��<G��<��<��<!��<o��<A��<���<f��<���<���<Ų�<���<���<f��<���<A��<t��<!��<`   `   ��<��<#��<L��<=��<��<��<#��<^��<���<^��<:��<���<���<X��<���<���<e��<���<���<E��<\��<���<h��<`   `   ұ�<
��<��<>��<��<
��<���<��<��<<��<S��<���<���<���<���<0��<���<���<Ͳ�<���<J��<<��<��<��<`   `   ��<��<���<��<��<���<��<Q��<?��<{��<���<���<���<V��<���<Ų�<f��<���<���<���<���<I��<N��<ܱ�<`   `   ��<��<G��<��<��<��<G��<��<|��<���<8��<E��<���<?��<��<?��<���<E��<J��<���<g��<��<Z��<��<`   `   ��<ñ�<ϱ�<��<��<��<��<��<?��<L��<^��<0��<}��<���<���<v��<A��<\��<<��<I��<��<ٱ�<��<��<`   `   ��<ұ�<���<߱�<ı�<��<V��<N��<��<���<���<e��<���<���<���<e��<t��<���<��<N��<Z��<��<���<߱�<`   `   ���<��<E��<��<��<��<��<"��<^��<��<��<g��<c��<]��<Z��<	��<!��<h��<��<ܱ�<��<��<߱�<9��<`   `   O��<i��<Q��<���<R��<���<���<���<Ҵ�<���<��<ɴ�<���<ɴ�<���<���<���<���<Ӵ�<���<0��<���<e��<i��<`   `   i��<���<\��<J��<���<���<t��<���<ݴ�<Ŵ�<���<���<���<���<���<��<ƴ�<c��<޴�<Ѵ�<Z��<O��<���<m��<`   `   Q��<\��<}��<V��<L��<A��<ڴ�<���<���<���<��<��<ش�<���<���<���<Դ�<A��<P��<V��<z��<\��<S��<���<`   `   ���<J��<V��<n��<}��<{��<���<���<���<c��<���<���<m��<���<���<{��<���<���<X��<I��<Z��<���<z��<���<`   `   R��<���<L��<}��<��<���<T��<Ҵ�<���<���<Ǵ�<���<���<Ҵ�<w��<���<���<}��<p��<���<=��<���<���<���<`   `   ���<���<A��<{��<���<���<���<���<���<���<���<���<���<���<w��<ȴ�<���<3��<޴�<���<(��<���<���<��<`   `   ���<t��<ڴ�<���<T��<���<��<z��<���<���<���<z��<��<���<T��<���<д�<t��<���<���<���<~��<Դ�<���<`   `   ���<���<���<���<Ҵ�<���<z��<���<״�<��<���<i��<���<��<���<���<ƴ�<���<޴�<ʴ�<s��<c��<Ĵ�<���<`   `   Ҵ�<ݴ�<���<���<���<���<���<״�<���<״�<���<���<���<���<���<ݴ�<���<���<��<���<ʹ�<���<o��<���<`   `   ���<Ŵ�<���<c��<���<���<���<��<״�<���<���<´�<m��<z��<���<´�<���<ٴ�<ٴ�<���<Ĵ�<��<Ӵ�<���<`   `   ��<���<��<���<Ǵ�<���<���<���<���<���<���<���<��<���<���<&��<���<��<д�<���<���<��<��<&��<`   `   ɴ�<���<��<���<���<���<z��<i��<���<´�<���<��<���<δ�<%��<ƴ�<ش�<ܴ�<��<���<��<���<���<8��<`   `   ���<���<ش�<m��<���<���<��<���<���<m��<��<���<y��<���<��<���<Y��<ϴ�<���<ϴ�<`��<���<s��<���<`   `   ɴ�<���<���<���<Ҵ�<���<���<��<���<z��<���<δ�<���<��<.��<(��<��<2��<��<���<7��<A��<��<���<`   `   ���<���<���<���<w��<w��<T��<���<���<���<���<%��<��<.��<8��<���<��<q��<��<���<��<.��<���<%��<`   `   ���<��<���<{��<���<ȴ�<���<���<ݴ�<´�<&��<ƴ�<���<(��<���<���<���<��<���<��<7��<���<���<%��<`   `   ���<ƴ�<Դ�<���<���<���<д�<ƴ�<���<���<���<ش�<Y��<��<��<���<���<���<��<��<S��<ش�<���<���<`   `   ���<c��<A��<���<}��<3��<t��<���<���<ٴ�<��<ܴ�<ϴ�<2��<q��<��<���<���<��<Ŵ�<��<��<Ӵ�<���<`   `   Ӵ�<޴�<P��<X��<p��<޴�<���<޴�<��<ٴ�<д�<��<���<��<��<���<��<��<���<��<���<ٴ�<z��<޴�<`   `   ���<Ѵ�<V��<I��<���<���<���<ʴ�<���<���<���<���<ϴ�<���<���<��<��<Ŵ�<��<���<Ĵ�<���<Ĵ�<���<`   `   0��<Z��<z��<Z��<=��<(��<���<s��<ʹ�<Ĵ�<���<��<`��<7��<��<7��<S��<��<���<Ĵ�<���<s��<ִ�<(��<`   `   ���<O��<\��<���<���<���<~��<c��<���<��<��<���<���<A��<.��<���<ش�<��<ٴ�<���<s��<m��<���<���<`   `   e��<���<S��<z��<���<���<Դ�<Ĵ�<o��<Ӵ�<��<���<s��<��<���<���<���<Ӵ�<z��<Ĵ�<ִ�<���<���<z��<`   `   i��<m��<���<���<���<��<���<���<���<���<&��<8��<���<���<%��<%��<���<���<޴�<���<(��<���<z��<��<`   `   ̶�<��<ж�<��<��<��<���<"��<���<c��<��<y��<���<y��<��<c��<t��<"��<,��<��<��<��<��<��<`   `   ��<��<ܶ�<ζ�<��<F��<���<��<?��<o��<���<F��<R��<���<X��<J��<��<��<+��<��<��<ζ�<߶�<��<`   `   ж�<ܶ�<L��<��<��<	��<���<���<��<��<���<-��<���<��<��<���<���<	��<��<��<G��<ܶ�<Ӷ�<ɶ�<`   `   ��<ζ�<��<m��<-��<��<#��<S��<V��<��<��<��<��<a��<=��<��<��<A��<S��<��<��<��<��<���<`   `   ��<��<��<-��<���<��<,��<G��<$��<M��<.��<M��<��<G��<T��<��<϶�<-��<
��<��<���<(��<���<(��<`   `   ��<F��<	��<��<��<}��<��<��<U��<4��<4��<`��<��<���<g��<)��<��<���<+��<��<��<���<��<���<`   `   ���<���<���<#��<,��<��<"��<.��<%��<߶�<��<.��<(��<��<.��<#��<��<���<��<��<N��<U��<i��<��<`   `   "��<��<���<S��<G��<��<.��<!��<��<��<!��<��<��<[��<=��<��<��<&��<>��<��<_��<L��<��<X��<`   `   ���<?��<��<V��<$��<U��<%��<��<ܶ�<��<7��<U��<��<V��<&��<?��<z��<o��<A��<���<���<���</��<o��<`   `   c��<o��<��<��<M��<4��<߶�<��<��<Ͷ�<4��<a��<��<q��<X��<h��<X��<^��<ڷ�<T��<g��<���<V��<<��<`   `   ��<���<���<��<.��<4��<��<!��<7��<4��<��<��<���<���<��<x��<`��<y��<˷�<���<���<y��<���<x��<`   `   y��<F��<-��<��<M��<`��<.��<��<U��<a��<��<��<R��<}��<���<Ʒ�<÷�<���<5��<O��<̷�<���<���<���<`   `   ���<R��<���<��<��<��<(��<��<��<��<���<R��<���<��<���<Է�<��<���<���<���<��<Է�<}��<��<`   `   y��<���<��<a��<G��<���<��<[��<V��<q��<���<}��<��<���<���<���<ŷ�<��<��<���<���<ַ�<��<ط�<`   `   ��<X��<��<=��<T��<g��<.��<=��<&��<X��<��<���<���<���<���<)��<��<!��<7��<)��<���<���<���<���<`   `   c��<J��<���<��<��<)��<#��<��<?��<h��<x��<Ʒ�<Է�<���<)��<D��<��<ɷ�<*��<?��<���<Ƿ�<���<x��<`   `   t��<��<���<��<϶�<��<��<��<{��<X��<`��<÷�<��<ŷ�<��<��<���<��<��<ŷ�<	��<÷�<h��<X��<`   `   "��<��<	��<A��<-��<���<���<&��<o��<^��<y��<���<���<��<!��<ɷ�<��<8��<��<���<̷�<y��<V��<{��<`   `   ,��<+��<��<S��<
��<+��<��<>��<A��<ڷ�<˷�<5��<���<��<7��<*��<��<��<۷�<5��<���<ڷ�<>��<>��<`   `   ��<��<��<��<��<��<��<��<���<T��<���<O��<���<���<)��<?��<ŷ�<���<5��<���<g��<���<��<���<`   `   ��<��<G��<��<���<��<N��<_��<���<g��<���<̷�<��<���<���<���<	��<̷�<���<g��<���<_��<i��<��<`   `   ��<ζ�<ܶ�<��<(��<���<U��<L��<���<���<y��<���<Է�<ַ�<���<Ƿ�<÷�<y��<ڷ�<���<_��<C��<��<;��<`   `   ��<߶�<Ӷ�<��<���<��<i��<��</��<V��<���<���<}��<��<���<���<h��<V��<>��<��<i��<��<���<��<`   `   ��<��<ɶ�<���<(��<���<��<X��<o��<<��<x��<���<��<ط�<���<x��<X��<{��<>��<���<��<;��<��<���<`   `   ��<a��<`��<J��<���<���<���<��<��<2��<ݹ�<F��<a��<F��<���<2��<���<��<ٹ�<���<���<J��<x��<a��<`   `   a��<N��<_��<O��<���<Թ�<��<���<��<Q��<��<��<��<��<9��<*��<���<ֹ�<���<���<d��<Q��<E��<f��<`   `   `��<_��<͹�<X��<L��<Ź�<J��<ӹ�<��<Թ�<��<ֹ�<���<Թ�<��<ӹ�<@��<Ź�<T��<X��<ǹ�<_��<e��<ֹ�<`   `   J��<O��<X��<ù�<ɹ�<���<���<��<��<߹�<��<��<��<���<���<���<���<޹�<���<I��<d��<N��<���<���<`   `   ���<���<L��<ɹ�<���<���<���<ɹ�<ٹ�<��<���<��<���<ɹ�<ù�<���<���<ɹ�<w��<���<���<���<D��<���<`   `   ���<Թ�<Ź�<���<���<��<���<���<۹�<���<���<��<���<���<��<Ϲ�<���<���<���<���<ع�<ɹ�<���<ù�<`   `   ���<��<J��<���<���<���<M��<ݹ�<��<	��<ֹ�<ݹ�<R��<���<���<���<;��<��<¹�<���<Թ�<���<��<���<`   `   ��<���<ӹ�<��<ɹ�<���<ݹ�<���< ��<��<���<ʹ�<���<ݹ�<���<Ź�<���<��<%��<߹�<���<���<ֹ�<B��<`   `   ��<��<��<��<ٹ�<۹�<��< ��<���< ��<���<۹�<���<��<��<��<���<'��<��<��</��<��<۹�<'��<`   `   2��<Q��<Թ�<߹�<��<���<	��<��< ��<���<���<'��<��<Ź�<9��<6��<-��<O��<W��<��<��<s��<F��<��<`   `   ݹ�<��<��<��<���<���<ֹ�<���<���<���<���<��<��<��<��<>��<d��<+��<R��<7��< ��<+��<���<>��<`   `   F��<��<ֹ�<��<��<��<ݹ�<ʹ�<۹�<'��<��<ǹ�<��<J��<?��<���<G��<��<s��<���<0��<)��<���<X��<`   `   a��<��<���<��<���<���<R��<���<���<��<��<��<O��<��<F��<���<���<���<j��<���<���<���<6��<��<`   `   F��<��<Թ�<���<ɹ�<���<���<ݹ�<��<Ź�<��<J��<��<K��<���<N��<���<���<ݺ�<l��<c��<Ѻ�<B��<���<`   `   ���<9��<��<���<ù�<��<���<���<��<9��<��<?��<F��<���<���<պ�<���<`��<���<պ�<_��<���<\��<?��<`   `   2��<*��<ӹ�<���<���<Ϲ�<���<Ź�<��<6��<>��<���<���<N��<պ�</��<���<v��<��<��<c��<���<���<?��<`   `   ���<���<@��<���<���<���<;��<���<���<-��<d��<G��<���<���<���<���<���<���<���<���<���<G��<l��<-��<`   `   ��<ֹ�<Ź�<޹�<ɹ�<���<��<��<'��<O��<+��<��<���<���<`��<v��<���<y��<ݺ�<x��<0��<+��<F��<2��<`   `   ٹ�<���<T��<���<w��<���<¹�<%��<��<W��<R��<s��<j��<ݺ�<���<��<���<ݺ�<���<s��<<��<W��<��<%��<`   `   ���<���<X��<I��<���<���<���<߹�<��<��<7��<���<���<l��<պ�<��<���<x��<s��<7��<��<��<ֹ�<���<`   `   ���<d��<ǹ�<d��<���<ع�<Թ�<���</��<��< ��<0��<���<c��<_��<c��<���<0��<<��<��<��<���<��<ع�<`   `   J��<Q��<_��<N��<���<ɹ�<���<���<��<s��<+��<)��<���<Ѻ�<���<���<G��<+��<W��<��<���<���<���<ƹ�<`   `   x��<E��<e��<���<D��<���<��<ֹ�<۹�<F��<���<���<6��<B��<\��<���<l��<F��<��<ֹ�<��<���<9��<���<`   `   a��<f��<ֹ�<���<���<ù�<���<B��<'��<��<>��<X��<��<���<?��<?��<-��<2��<%��<���<ع�<ƹ�<���<ǹ�<`   `   ��<ݻ�<ܻ�<���<4��<<��<K��<���<���<Ӽ�<��<9��<
��<9��<��<Ӽ�<���<���<{��<<��<��<���<���<ݻ�<`   `   ݻ�<!��<+��<��<���<���<c��<\��<Ǽ�<��<ڼ�<޼�<��<ڼ�<׼�<Ҽ�<z��<P��<}��<���<!��<��<��<��<`   `   ܻ�<+��<9��<"��< ��<	��<���<}��<m��<^��<��<��<޼�<^��<z��<}��<���<	��<)��<"��<3��<+��<��<���<`   `   ���<��<"��<y��<E��<��<T��<˼�<���<~��<���<���<���<���<���<A��<1��<Z��<\��<��<!��<��<���<��<`   `   4��<���< ��<E��<���<���<1��<���<���<���<_��<���<���<���<]��<���<���<E��<L��<���<��<��<8��<��<`   `   <��<���<	��<��<���<~��<V��<i��<v��<���<���<���<w��<C��<e��<μ�<1��<���<}��<@��<��<e��<\��<ֻ�<`   `   K��<c��<���<T��<1��<V��<ʼ�<5��<n��<���<c��<5��<м�<V��<6��<T��<���<c��<d��<Y��<���<S��<���<Y��<`   `   ���<\��<}��<˼�<���<i��<5��<=��<`��<k��<<��<"��<w��<���<���<n��<z��<���<ּ�<��<˼�<���<���<��<`   `   ���<Ǽ�<m��<���<���<v��<n��<`��<��<`��<���<v��<{��<���<���<Ǽ�<���<���<l��<ڼ�</��<ڼ�<X��<���<`   `   Ӽ�<��<^��<~��<���<���<���<k��<`��<y��<���<���<���<O��<׼�<׼�<���<��<���<��<��<��<��<���<`   `   ��<ڼ�<��<���<_��<���<c��<<��<���<���<K��<���<��<ڼ�<���<��<G��<x��<���<���<X��<x��<n��<��<`   `   9��<޼�<��<���<���<���<5��<"��<v��<���<���<��<��<=��<���<!��<+��<���<u��<���<���<��<��<���<`   `   
��<��<޼�<���<���<w��<м�<w��<{��<���<��<��<���<,��<A��<6��<(��<˽�<��<˽�<1��<6��<1��<,��<`   `   9��<ڼ�<^��<���<���<C��<V��<���<���<O��<ڼ�<=��<,��<k��<Ľ�<���<ǽ�<$��<��<���<���<ݽ�<b��<��<`   `   ��<׼�<z��<���<]��<e��<6��<���<���<׼�<���<���<A��<Ľ�<��<���<���<J��<��<���<���<Ľ�<X��<���<`   `   Ӽ�<Ҽ�<}��<A��<���<μ�<T��<n��<Ǽ�<׼�<��<!��<6��<���<���<���<��<��<ܽ�<ǽ�<���<(��<��<��<`   `   ���<z��<���<1��<���<1��<���<z��<���<���<G��<+��<(��<ǽ�<���<��<s��<��<���<ǽ�<!��<+��<O��<���<`   `   ���<P��<	��<Z��<E��<���<c��<���<���<��<x��<���<˽�<$��<J��<��<��<b��<��<���<���<x��<��<���<`   `   {��<}��<)��<\��<L��<}��<d��<ּ�<l��<���<���<u��<��<��<��<ܽ�<���<��<D��<u��<t��<���<i��<ּ�<`   `   <��<���<"��<��<���<@��<Y��<��<ڼ�<��<���<���<˽�<���<���<ǽ�<ǽ�<���<u��<���<��<��<���<F��<`   `   ��<!��<3��<!��<��<��<���<˼�</��<��<X��<���<1��<���<���<���<!��<���<t��<��<��<˼�<���<��<`   `   ���<��<+��<��<��<e��<S��<���<ڼ�<��<x��<��<6��<ݽ�<Ľ�<(��<+��<x��<���<��<˼�<@��<\��<3��<`   `   ���<��<��<���<8��<\��<���<���<X��<��<n��<��<1��<b��<X��<��<O��<��<i��<���<���<\��<-��<���<`   `   ݻ�<��<���<��<��<ֻ�<Y��<��<���<���<��<���<,��<��<���<��<���<���<ּ�<F��<��<3��<���<���<`   `   ���<l��<���<ؾ�<׾�<��<��<���<��<ѿ�<w��<���<��<���<���<ѿ�<ۿ�<���<��<��<���<ؾ�<���<l��<`   `   l��<g��<Y��<T��<���<��<��<5��<���<��<���<���<���<���<̿�<���<Q��<
��<��<ž�<h��<K��<_��<p��<`   `   ���<Y��<���<���<���<(��<���<<��<A��<Կ�<��<[��<ֿ�<Կ�<M��<<��<���<(��<���<���<���<Y��<���<S��<`   `   ؾ�<T��<���<,��<��<��<6��<p��<t��<e��<*��<*��<r��<��<Y��<#��<	��<(��<��<���<h��<ܾ�<ľ�<̾�<`   `   ׾�<���<���<��<پ�<
��<��<U��<*��<Z��<\��<Z��<��<U��</��<
��<���<��<̾�<���<���<־�<���<־�<`   `   ��<��<(��<��<
��<V��<0��<��<^��<p��<p��<i��<)��<��<?��<��<	��<��<��<#��<
��<	��<��<���<`   `   ��<��<���<6��<��<0��<M��<>��<S��<���<H��<>��<S��<0��<��<6��<���<��< ��<��<>��<��<Z��<��<`   `   ���<5��<<��<p��<U��<��<>��<���<I��<T��<���<+��<)��<i��<Y��<-��<Q��<���<Z��<p��<;��<'��<g��<u��<`   `   ��<���<A��<t��<*��<^��<S��<I��<F��<I��<f��<^��<	��<t��<g��<���<��<ܿ�<���<ο�<���<ο�<y��<ܿ�<`   `   ѿ�<��<Կ�<e��<Z��<p��<���<T��<I��<���<p��<n��<r��<ƿ�<̿�<տ�<ؿ�<$��<��<���<���<-��<��<���<`   `   w��<���<��<*��<\��<p��<H��<���<f��<p��<I��<*��<��<���<���<޿�<.��<��<��<=��<ٿ�<��<R��<޿�<`   `   ���<���<[��<*��<Z��<i��<>��<+��<^��<n��<*��<L��<���<���<$��<c��<6��<��<���<���<��<��<[��<;��<`   `   ��<���<ֿ�<r��<��<)��<S��<)��<	��<r��<��<���<��<C��<o��<x��<���<���<���<���<���<x��<`��<C��<`   `   ���<���<Կ�<��<U��<��<0��<i��<t��<ƿ�<���<���<C��<���<U��<���<t��<���<���<X��<���<l��<z��<6��<`   `   ���<̿�<M��<Y��</��<?��<��<Y��<g��<̿�<���<$��<o��<U��<���<'��<���<A��<���<'��<���<U��<���<$��<`   `   ѿ�<���<<��<#��<
��<��<5��<-��<���<տ�<޿�<c��<x��<���<'��<}��<���<���<c��<>��<���<k��<[��<߿�<`   `   ۿ�<Q��<���<	��<���<	��<���<Q��<��<ؿ�<.��<6��<���<t��<���<���<���<���<���<t��<���<6��<6��<ؿ�<`   `   ���<
��<(��<(��<��<��<��<���<ܿ�<$��<��<��<���<���<A��<���<���<X��<���<���<��<��<��<��<`   `   ��<��<���<��<̾�<��< ��<Z��<���<��<��<���<���<���<���<c��<���<���<���<���<���<��<���<Z��<`   `   ��<ž�<���<���<���<#��<��<p��<ο�<���<=��<���<���<X��<'��<>��<t��<���<���<=��<���<ڿ�<g��<
��<`   `   ���<h��<���<h��<���<
��<>��<;��<���<���<ٿ�<��<���<���<���<���<���<��<���<���<���<;��<Y��<
��<`   `   ؾ�<K��<Y��<ܾ�<־�<	��<��<'��<ο�<-��<��<��<x��<l��<U��<k��<6��<��<��<ڿ�<;��<��<��<��<`   `   ���<_��<���<ľ�<���<��<Z��<g��<y��<��<R��<[��<`��<z��<���<[��<6��<��<���<g��<Y��<��<t��<ľ�<`   `   l��<p��<S��<̾�<־�<���<��<u��<ܿ�<���<޿�<;��<C��<6��<$��<߿�<ؿ�<��<Z��<
��<
��<��<ľ�<D��<`   `   ���<���<��<2��<a��<���<���<8��<r��<���<���<��<���<��<��<���<O��<8��<��<���<>��<2��<,��<���<`   `   ���<��<���<I��<Z��<���<���<���<D��<���<���<���<���<���<���<O��<���<���<���<l��<Z��<���<���<���<`   `   ��<���<
��<���<3��<���<#��<)��<��<6��<���<s��<|��<6��<"��<)��<��<���<8��<���<��<���<��<���<`   `   2��<I��<���<z��<���<���<���<5��<��<2��<���<���<<��<"��<"��<���<���<���<c��<���<Z��<7��<��<��<`   `   a��<Z��<3��<���<���<���<���<��< ��<#��<E��<#��<���<��<���<���<���<���<X��<Z��<L��<A��<���<A��<`   `   ���<���<���<���<���<;��<���<��<��<��<��<��<��<���<(��<
��<���<���<���<���<���<���<���<���<`   `   ���<���<#��<���<���<���<��<���<���<���<���<���<��<���<���<���<��<���<���<���< ��<��<��<���<`   `   8��<���<)��<5��<��<��<���<���<���<���<���<���<��<!��<"��<��<���<=��<L��<,��<7��<&��<&��<c��<`   `   r��<D��<��<��< ��<��<���<���<���<���<���<��<���<��<:��<D��<U��<��<p��<���<���<���<`��<��<`   `   ���<���<6��<2��<#��<��<���<���<���<���<��<5��<<��<(��<���<���<v��<���<L��<	��<��<c��<���<_��<`   `   ���<���<���<���<E��<��<���<���<���<��<2��<���<���<���<��<2��<,��<a��<���<n��<[��<a��<J��<2��<`   `   ��<���<s��<���<#��<��<���<���<��<5��<���<e��<���<��<"��<���<���<���<���<���<���<���<���<5��<`   `   ���<���<|��<<��<���<��<��<��<���<<��<���<���<}��< ��<c��<���<M��<"��<%��<"��<U��<���<V��< ��<`   `   ��<���<6��<"��<��<���<���<!��<��<(��<���<��< ��<���<��<��<E��<���<���<.��<$��<��<���<���<`   `   ��<���<"��<"��<���<(��<���<"��<:��<���<��<"��<c��<��<%��<{��<8��<���<g��<{��<��<��<s��<"��<`   `   ���<O��<)��<���<���<
��<���<��<D��<���<2��<���<���<��<{��<���<���<���<z��<���<$��<���<���<1��<`   `   O��<���<��<���<���<���<��<���<U��<v��<,��<���<M��<E��<8��<���<��<���<<��<E��<G��<���<3��<v��<`   `   8��<���<���<���<���<���<���<=��<��<���<a��<���<"��<���<���<���<���<���<���<��<���<`��<���<���<`   `   ��<���<8��<c��<X��<���<���<L��<p��<L��<���<���<%��<���<g��<z��<<��<���<F��<���<s��<L��<l��<L��<`   `   ���<l��<���<���<Z��<���<���<,��<���<	��<n��<���<"��<.��<{��<���<E��<��<���<n��<��<���<&��<���<`   `   >��<Z��<��<Z��<L��<���< ��<7��<���<��<[��<���<U��<$��<��<$��<G��<���<s��<��<���<7��<��<���<`   `   2��<���<���<7��<A��<���<��<&��<���<c��<a��<���<���<��<��<���<���<`��<L��<���<7��<���<���<S��<`   `   ,��<���<��<��<���<���<��<&��<`��<���<J��<���<V��<���<s��<���<3��<���<l��<&��<��<���<���<��<`   `   ���<���<���<��<A��<���<���<c��<��<_��<2��<5��< ��<���<"��<1��<v��<���<L��<���<���<S��<��<���<`   `   ��<w��<p��<���<
��<0��<���<A��<���<���<���<1��<,��<1��<��<���<~��<A��<���<0��<���<���<���<w��<`   `   w��<���<J��<���<D��<���<���<!��<r��<���<���<���<���<���<���<|��<2��<���<���<T��<���<=��<���<}��<`   `   p��<J��<���<���<+��<f��<���<;��<4��<F��<z��<T��<u��<F��<8��<;��<���<f��<,��<���<���<J��<n��<4��<`   `   ���<���<���<��<z��</��<���<��</��<?��<D��<B��<E��<9��<��<���<A��<���<
��<���<���<���<���<���<`   `   
��<D��<+��<z��<���<���<���<���<��<���<���<���<���<���<���<���<���<z��<H��<D��<���<,��<<��<,��<`   `   0��<���<f��</��<���<���<q��<���<���<���<���<���<���<b��<���<���<A��<Z��<���<5��<���<O��<L��<���<`   `   ���<���<���<���<���<q��<���<���<��<8��<���<���<��<q��<��<���<���<���<���<���<���<���<���<���<`   `   A��<!��<;��<��<���<���<���<���<���<���<���<���<���<���<��<.��<2��<G��<\��<[��<;��</��<W��<l��<`   `   ���<r��<4��</��<��<���<��<���<>��<���<��<���<���</��<O��<r��<���<���<j��<���<���<���<]��<���<`   `   ���<���<F��<?��<���<���<8��<���<���<)��<���<���<E��<:��<���<���<���<��<���<���<���<��<��<���<`   `   ���<���<z��<D��<���<���<���<���<��<���<���<D��<���<���<���<4��<���<���<���<���<���<���<���<4��<`   `   1��<���<T��<B��<���<���<���<���<���<���<D��<G��<���<7��<x��<}��<���<��<���<��< ��<���<z��<���<`   `   ,��<���<u��<E��<���<���<��<���<���<E��<���<���< ��<x��<���<���<]��<W��<���<W��<c��<���<���<x��<`   `   1��<���<F��<9��<���<b��<q��<���</��<:��<���<7��<x��<A��<s��<D��<���<���<���<���<P��<���<=��<r��<`   `   ��<���<8��<��<���<���<��<��<O��<���<���<x��<���<s��<i��<���<��< ��<$��<���<O��<s��<���<x��<`   `   ���<|��<;��<���<���<���<���<.��<r��<���<4��<}��<���<D��<���<"��<��<��<��<���<P��<���<z��<2��<`   `   ~��<2��<���<A��<���<A��<���<2��<���<���<���<���<]��<���<��<��<���<��<��<���<Y��<���<���<���<`   `   A��<���<f��<���<z��<Z��<���<G��<���<��<���<��<W��<���< ��<��<��<.��<���<P��< ��<���<��<���<`   `   ���<���<,��<
��<H��<���<���<\��<j��<���<���<���<���<���<$��<��<��<���<���<���<���<���<c��<\��<`   `   0��<T��<���<���<D��<5��<���<[��<���<���<���<��<W��<���<���<���<���<P��<���<���<���<���<W��<w��<`   `   ���<���<���<���<���<���<���<;��<���<���<���< ��<c��<P��<O��<P��<Y��< ��<���<���<���<;��<���<���<`   `   ���<=��<J��<���<,��<O��<���</��<���<��<���<���<���<���<s��<���<���<���<���<���<;��<���<L��<<��<`   `   ���<���<n��<���<<��<L��<���<W��<]��<��<���<z��<���<=��<���<z��<���<��<c��<W��<���<L��<0��<���<`   `   w��<}��<4��<���<,��<���<���<l��<���<���<4��<���<x��<r��<x��<2��<���<���<\��<w��<���<<��<���<(��<`   `   j��<���<���<'��<���<��<g��<���<`��<���<���<U��<F��<U��<���<���<M��<���<}��<��<���<'��<���<���<`   `   ���<���<(��<U��<���<��<���<���<<��<���<
��<��<��<��<���<E��<���<���<��<���<\��<��<���<���<`   `   ���<(��<c��<q��<���<��<���<x��<���<r��<���<���<���<r��<���<x��<���<��<���<q��<g��<(��<���<���<`   `   '��<U��<q��<���<���<6��<���<���<���<���<��<��<��<���<���<���<@��<���<���<g��<\��<-��<���<���<`   `   ���<���<���<���<���<M��<���<���<���<(��<'��<(��<���<���<���<M��<���<���<���<���<���<s��<'��<s��<`   `   ��<��<��<6��<M��<|��<���<L��<���<���<���<���<O��<���<u��<Z��<@��<��<��<��<��<���<���<��<`   `   g��<���<���<���<���<���<���<l��<Z��<��<N��<l��<���<���<���<���<���<���<k��<���<���<L��<���<���<`   `   ���<���<x��<���<���<L��<l��<���<j��<s��<���<`��<O��<���<���<n��<���<���<���<2��<���<���<1��<���<`   `   `��<<��<���<���<���<���<Z��<j��<���<j��<c��<���<���<���<���<<��<P��<{��<���<���<��<���<���<{��<`   `   ���<���<r��<���<(��<���<��<s��<j��<���<���<5��<��<h��<���<���<6��<u��<x��<���<���<���<t��<,��<`   `   ���<
��<���<��<'��<���<N��<���<c��<���<��<��<���<
��<���<V��<���<���<��<<��<���<���<���<V��<`   `   U��<��<���<��<(��<���<l��<`��<���<5��<��<���<��<[��<���<d��<}��<���< ��<*��<���<r��<c��<���<`   `   F��<��<���<��<���<O��<���<O��<���<��<���<��<=��<���<���<"��<f��<u��<���<u��<j��<"��<���<���<`   `   U��<��<r��<���<���<���<���<���<���<h��<
��<[��<���<"��<���<���<���<���<���<���<���<���<"��<���<`   `   ���<���<���<���<���<u��<���<���<���<���<���<���<���<���<���<��<��<:��<,��<��<���<���<���<���<`   `   ���<E��<x��<���<M��<Z��<���<n��<<��<���<V��<d��<"��<���<��<���<_��<U��<���<��<���<��<c��<S��<`   `   M��<���<���<@��<���<@��<���<���<P��<6��<���<}��<f��<���<��<_��<l��<_��<��<���<c��<}��<���<6��<`   `   ���<���<��<���<���<��<���<���<{��<u��<���<���<u��<���<:��<U��<_��<B��<���<r��<���<���<t��<���<`   `   }��<��<���<���<���<��<k��<���<���<x��<��< ��<���<���<,��<���<��<���<���< ��<
��<x��<���<���<`   `   ��<���<q��<g��<���<��<���<2��<���<���<<��<*��<u��<���<��<��<���<r��< ��<9��<���<���<1��<���<`   `   ���<\��<g��<\��<���<��<���<���<��<���<���<���<j��<���<���<���<c��<���<
��<���<���<���<���<��<`   `   '��<��<(��<-��<s��<���<L��<���<���<���<���<r��<"��<���<���<��<}��<���<x��<���<���<?��<���<���<`   `   ���<���<���<���<'��<���<���<1��<���<t��<���<c��<���<"��<���<c��<���<t��<���<1��<���<���<��<���<`   `   ���<���<���<���<s��<��<���<���<{��<,��<V��<���<���<���<���<S��<6��<���<���<���<��<���<���<���<`   `   ���<���<���<U��<���<���<���<��<���<n��<z��<���<���<���<��<n��<���<��<���<���<���<U��<��<���<`   `   ���<~��<2��<t��<��<���<R��<���<���<���<���<>��<=��<���<���<���<���<J��<���<��<t��<+��<���<���<`   `   ���<2��<��<���<:��<���<^��<���<J��<6��<n��<���<s��<6��<D��<���<d��<���<3��<���<���<2��<���<]��<`   `   U��<t��<���<Q��<~��<'��<U��<���<��<���<���<���<���<$��<���<M��<)��<���<O��<���<t��<Z��<x��<u��<`   `   ���<��<:��<~��<���<���<<��<���<���<���<���<���<���<���<E��<���<���<~��<C��<��<���<���<���<���<`   `   ���<���<���<'��<���<���<Q��<?��<���<t��<x��<���<>��<H��<���<��<)��<���<���<���<s��<���<���<s��<`   `   ���<R��<^��<U��<<��<Q��<n��<h��<u��<B��<j��<h��<x��<Q��<4��<U��<d��<R��<���<��<?��<���<=��<��<`   `   ��<���<���<���<���<?��<h��<[��<]��<d��<_��<`��<>��<���<���<���<���<$��<"��<���<��<��<���<$��<`   `   ���<���<J��<��<���<���<u��<]��<@��<]��<z��<���<���<��<R��<���<���<���<��<��<���<��<���<���<`   `   n��<���<6��<���<���<t��<B��<d��<]��<:��<x��<��<���<.��<���<s��<c��<���<(��<���<���<*��<���<a��<`   `   z��<���<n��<���<���<x��<j��<_��<z��<x��<���<���<v��<���<v��<���<9��<���<���<���<���<���<9��<���<`   `   ���<>��<���<���<���<���<h��<`��<���<��<���<���<=��<���<n��<���<=��<���<���<���<���<;��<���<o��<`   `   ���<=��<s��<���<���<>��<x��<>��<���<���<v��<=��<���<���<���<���<��<7��<e��<7��<��<���<���<���<`   `   ���<���<6��<$��<���<H��<Q��<���<��<.��<���<���<���</��<���<{��<���<��<��<���<|��<���<2��<���<`   `   ��<���<D��<���<E��<���<4��<���<R��<���<v��<n��<���<���<���<���<O��<���<S��<���<���<���<���<n��<`   `   n��<���<���<M��<���<��<U��<���<���<s��<���<���<���<{��<���<f��<���<���<d��<���<|��<���<���<���<`   `   ���<���<d��<)��<���<)��<d��<���<���<c��<9��<=��<��<���<O��<���<��<���<P��<���<��<=��<;��<c��<`   `   ��<J��<���<���<~��<���<R��<$��<���<���<���<���<7��<��<���<���<���<���<��<8��<���<���<���<���<`   `   ���<���<3��<O��<C��<���<���<"��<��<(��<���<���<e��<��<S��<d��<P��<��<e��<���<���<(��<���<"��<`   `   ���<��<���<���<��<���<��<���<��<���<���<���<7��<���<���<���<���<8��<���<���<���<��<���<��<`   `   ���<t��<���<t��<���<s��<?��<��<���<���<���<���<��<|��<���<|��<��<���<���<���<���<��<E��<s��<`   `   U��<+��<2��<Z��<���<���<���<��<��<*��<���<;��<���<���<���<���<=��<���<(��<��<��<���<���<���<`   `   ��<���<���<x��<���<���<=��<���<���<���<9��<���<���<2��<���<���<;��<���<���<���<E��<���<���<x��<`   `   ���<���<]��<u��<���<s��<��<$��<���<a��<���<o��<���<���<n��<���<c��<���<"��<��<s��<���<x��<U��<`   `   G��<���<���<���<[��<��<���<���<���<A��<$��<���<6��<���<#��<A��<���<���<���<��<]��<���<���<���<`   `   ���<���<O��<���<���<G��<���<���<T��<���<���<���<���<���<���<X��<���<���<M��<���<���<L��<���<���<`   `   ���<O��<a��<	��<���<Y��<���<���<(��<���<	��<���<��<���<��<���<���<Y��<���<	��<j��<O��<���<���<`   `   ���<���<	��<j��<���<���<���<R��<���<<��<���<���<7��<���<X��<���<���<���<p��<��<���<���<$��<��<`   `   [��<���<���<���<U��<���<���<��<f��<���<���<���<g��<��<���<���<W��<���<���<���<\��<X��<��<X��<`   `   ��<G��<Y��<���<���<'��<��</��<4��<��<��<7��<*��<��<-��<���<���<U��<M��<��<��<���<���<��<`   `   ���<���<���<���<���<��<��<���<��<���<��<���<��<��<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<R��<��</��<���<w��<���<���<|��<���<*��<��<X��<���<���<���<-��<6��<i��<n��<;��<'��<`   `   ���<T��<(��<���<f��<4��<��<���<@��<���<��<4��<h��<���<&��<T��<���<��<O��<:��<R��<:��<P��<��<`   `   A��<���<���<<��<���<��<���<���<���<���<��<���<7��<���<���<F��<���<��<K��<���<���<E��<��<���<`   `   $��<���<	��<���<���<��<��<|��<��<��<}��<���<��<���<��<���<]��<���<��<,��<��<���<R��<���<`   `   ���<���<���<���<���<7��<���<���<4��<���<���<���<���<���<��<���<���<���<!��<��<���<���<���<��<`   `   6��<���<��<7��<g��<*��<��<*��<h��<7��<��<���<6��<`��<7��<���<���<���<���<���<��<���<8��<`��<`   `   ���<���<���<���<��<��<��<��<���<���<���<���<`��<���<���<��<��<���<���<��<��<���<���<f��<`   `   #��<���<��<X��<���<-��<���<X��<&��<���<��<��<7��<���<��<��<���<D��<���<��<)��<���<-��<��<`   `   A��<X��<���<���<���<���<���<���<T��<F��<���<���<���<��<��<���<���<���<���<��<��<���<���<���<`   `   ���<���<���<���<W��<���<���<���<���<���<]��<���<���<��<���<���<��<���<���<��<���<���<]��<���<`   `   ���<���<Y��<���<���<U��<���<���<��<��<���<���<���<���<D��<���<���<>��<���<���<���<���<��< ��<`   `   ���<M��<���<p��<���<M��<���<-��<O��<K��<��<!��<���<���<���<���<���<���<���<!��<��<K��<F��<-��<`   `   ��<���<	��<��<���<��<���<6��<:��<���<,��<��<���<��<��<��<��<���<!��<(��<���<>��<;��<���<`   `   ]��<���<j��<���<\��<��<���<i��<R��<���<��<���<��<��<)��<��<���<���<��<���<S��<i��<���<��<`   `   ���<L��<O��<���<X��<���<���<n��<:��<E��<���<���<���<���<���<���<���<���<K��<>��<i��<���<���<\��<`   `   ���<���<���<$��<��<���<���<;��<P��<��<R��<���<8��<���<-��<���<]��<��<F��<;��<���<���<��<$��<`   `   ���<���<���<��<X��<��<���<'��<��<���<���<��<`��<f��<��<���<���< ��<-��<���<��<\��<$��<���<`   `   ���<��<���<#��<���<R��<���<���<��<��<���<W��<���<W��<���<��<��<���<���<R��<���<#��<���<��<`   `   ��<I��<���<���<C��<h��<���<���<���<b��<��<@��<8��<	��<m��<���<���<���<u��<@��<���<���<P��<!��<`   `   ���<���<u��<!��<���<���<���<���<C��<���<���<���<���<���<7��<���<���<���<���<!��<��<���<���<���<`   `   #��<���<!��<u��<h��<	��<���<.��<���<���<��<��<���<���<:��<���<���<e��<���<"��<���<&��<��<��<`   `   ���<C��<���<h��<���<��<���<-��<O��<���<��<���<X��<-��<���<��<���<h��<���<C��<���<���<5��<���<`   `   R��<h��<���<	��<��<���<���<$��<��<��<��<��<��<���<���<��<���<���<u��<U��<c��<&��<-��<m��<`   `   ���<���<���<���<���<���<u��<���<���<���<���<���<{��<���<���<���<���<���<���<���<���<Q��<���<���<`   `   ���<���<���<.��<-��<$��<���<���<���<���<���<���<��<+��<:��<���<���<���<���<��<��<��<"��<���<`   `   ��<���<C��<���<O��<��<���<���<���<���<���<��<[��<���<6��<���<��<k��<���<���<���<���<���<k��<`   `   ��<b��<���<���<���<��<���<���<���<���<��<���<���<���<m��<��<���<��<\��<���<���<N��<&��<���<`   `   ���<��<���<��<��<��<���<���<���<��<��<��<���<��<���<v��<��<���<���<��<���<���<��<v��<`   `   W��<@��<���<��<���<��<���<���<��<���<��<���<8��<Z��<��<2��<���<D��<���<���<9��<���<8��<��<`   `   ���<8��<���<���<X��<��<{��<��<[��<���<���<8��<���<���<���<��<9��<���<e��<���<6��<��<���<���<`   `   W��<	��<���<���<-��<���<���<+��<���<���<��<Z��<���<���<���<��<���<���<���<���<��<���<���<���<`   `   ���<m��<7��<:��<���<���<���<:��<6��<m��<���<��<���<���<��<"��<���<���<���<"��</��<���<���<��<`   `   ��<���<���<���<��<��<���<���<���<��<v��<2��<��<��<"��<���<���<���<���<��<��<
��<8��<r��<`   `   ��<���<���<���<���<���<���<���<��<���<��<���<9��<���<���<���<���<���<���<���<;��<���<��<���<`   `   ���<���<���<e��<h��<���<���<���<k��<��<���<D��<���<���<���<���<���<���<���<���<9��<���<&��<k��<`   `   ���<u��<���<���<���<u��<���<���<���<\��<���<���<e��<���<���<���<���<���<O��<���<���<\��<���<���<`   `   R��<@��<!��<"��<C��<U��<���<��<���<���<��<���<���<���<"��<��<���<���<���<��<���<���<"��<���<`   `   ���<���<��<���<���<c��<���<��<���<���<���<9��<6��<��</��<��<;��<9��<���<���<���<��<���<c��<`   `   #��<���<���<&��<���<&��<Q��<��<���<N��<���<���<��<���<���<
��<���<���<\��<���<��<S��<-��<���<`   `   ���<P��<���<��<5��<-��<���<"��<���<&��<��<8��<���<���<���<8��<��<&��<���<"��<���<-��<0��<��<`   `   ��<!��<���<��<���<m��<���<���<k��<���<v��<��<���<���<��<r��<���<k��<���<���<c��<���<��<���<`   `   ���<���<���<���<���<���<w��<���<��<���<���<��<���<��<���<���<7��<���<[��<���<���<���<���<���<`   `   ���<���<���<R��<S��<���<'��<h��<���<���<��<��<��<��<���<���<T��<0��<���<J��<D��<���<���<���<`   `   ���<���<���<���<���<���<���<��<G��<��<���<��<���<��<;��<��<���<���<���<���<���<���<���<d��<`   `   ���<R��<���<f��<y��<|��<J��<���<���<M��<G��<D��<C��<���<���<S��<h��<o��<y��<���<D��<���<T��<L��<`   `   ���<S��<���<y��<���<���<F��<���<
��<!��<h��<!��<��<���<,��<���<��<y��<���<S��<���<s��<���<s��<`   `   ���<���<���<|��<���<���<��<���<u��<���<���<q��<w��<'��<���<��<h��<���<���<���<��<I��<Q��<,��<`   `   w��<'��<���<J��<F��<��<���<,��<'��<���<)��<,��<���<��<>��<J��<���<'��<d��<���<��<e��<���<���<`   `   ���<h��<��<���<���<���<,��<b��<���<���<e��<4��<w��<���<���<��<T��<���<���<���<4��<C��<���<���<`   `   ��<���<G��<���<
��<u��<'��<���<���<���<��<u��<��<���<0��<���<2��<���<H��<W��<5��<W��<T��<���<`   `   ���<���<��<M��<!��<���<���<���<���<���<���<��<C��<��<���<���<a��<+��<���<���<���<���<2��<u��<`   `   ���<��<���<G��<h��<���<)��<e��<��<���<o��<G��<���<��<���<���<���<���<���<���<��<���<r��<���<`   `   ��<��<��<D��<!��<q��<,��<4��<u��<��<G��<��<��<��<���<���<��<��<��<���<��<��<���<���<`   `   ���<��<���<C��<��<w��<���<w��<��<C��<���<��<���<c��<���<��<���<���<F��<���<���<��<��<c��<`   `   ��<��<��<���<���<'��<��<���<���<��<��<��<c��<���<���<E��<���<S��<f��<���<7��<v��<���<n��<`   `   ���<���<;��<���<,��<���<>��<���<0��<���<���<���<���<���<���<���<���<%��<_��<���<���<���<���<���<`   `   ���<���<��<S��<���<��<J��<��<���<���<���<���<��<E��<���<q��<F��<Z��<���<���<7��<(��<���<���<`   `   7��<T��<���<h��<��<h��<���<T��<2��<a��<���<��<���<���<���<F��<���<F��<���<���<���<��<���<a��<`   `   ���<0��<���<o��<y��<���<'��<���<���<+��<���<��<���<S��<%��<Z��<F��<��<f��< ��<��<���<2��<���<`   `   [��<���<���<y��<���<���<d��<���<H��<���<���<��<F��<f��<_��<���<���<f��<(��<��<���<���<D��<���<`   `   ���<J��<���<���<S��<���<���<���<W��<���<���<���<���<���<���<���<���< ��<��<���<���<R��<���<��<`   `   ���<D��<���<D��<���<��<��<4��<5��<���<��<��<���<7��<���<7��<���<��<���<���<H��<4��<��<��<`   `   ���<���<���<���<s��<I��<e��<C��<W��<���<���<��<��<v��<���<(��<��<���<���<R��<4��<m��<Q��<i��<`   `   ���<���<���<T��<���<Q��<���<���<T��<2��<r��<���<��<���<���<���<���<2��<D��<���<��<Q��<���<T��<`   `   ���<���<d��<L��<s��<,��<���<���<���<u��<���<���<c��<n��<���<���<a��<���<���<��<��<i��<T��<k��<`   `   ��<���<���<8��<��<��<+��<���<���<^��<a��<���<���<���<N��<^��<���<���<��<��<1��<8��<���<���<`   `   ���<���<���<���<o��<)��<V��<���<���<6��<f��<���<���<e��<K��<���<���<e��<A��<^��<���<���<���<���<`   `   ���<���< ��<���<���<���<?��<?��<e��<��<���<���<���<��<Y��<?��<H��<���<���<���<��<���<���<[��<`   `   8��<���<���<���<���<g��<���<T��<B��<:��<5��<4��<.��<9��<h��<���<N��<���<���<���<���<5��<���<���<`   `   ��<o��<���<���<���<���<}��<���<���<���<���<���<���<���<Y��<���<���<���<o��<o��<$��<���<���<���<`   `   ��<)��<���<g��<���<��<���<���<��<^��<_��<���<���<���< ��<���<N��<��<A��<��< ��<���<���<��<`   `   +��<V��<?��<���<}��<���<���<Z��<���<���<���<Z��<���<���<y��<���<L��<V��<��<C��<'��<B��<��<C��<`   `   ���<���<?��<T��<���<���<Z��<T��<M��<D��<T��<i��<���<���<h��<K��<���<���<���<i��<i��<{��<p��<���<`   `   ���<���<e��<B��<���<��<���<M��<W��<M��<���<��<���<B��<E��<���<���<T��<��<;��<��<;��< ��<T��<`   `   ^��<6��<��<:��<���<^��<���<D��<M��<���<_��<���<.��<(��<K��<[��<���<&��<{��<��<n��<c��<.��<���<`   `   a��<f��<���<5��<���<_��<���<T��<���<_��<���<5��<���<f��<P��<u��<���<o��<��<���<F��<o��<���<u��<`   `   ���<���<���<4��<���<���<Z��<i��<��<���<5��<��<���<���<���<;��<���<���<���<���<���<���<C��<���<`   `   ���<���<���<.��<���<���<���<���<���<.��<���<���<���<;��<q��<��<8��<l��<���<l��<1��<��<~��<;��<`   `   ���<e��<��<9��<���<���<���<���<B��<(��<f��<���<;��<���<���<���<��<B��<Z��<7��<���<���<���<F��<`   `   N��<K��<Y��<h��<Y��< ��<y��<h��<E��<K��<P��<���<q��<���<���<���<���<���<���<���<���<���<^��<���<`   `   ^��<���<?��<���<���<���<���<K��<���<[��<u��<;��<��<���<���<��<2��<K��<-��<p��<���<��<C��<u��<`   `   ���<���<H��<N��<���<N��<L��<���<���<���<���<���<8��<��<���<2��<��<2��<���<��<>��<���<���<���<`   `   ���<e��<���<���<���<��<V��<���<T��<&��<o��<���<l��<B��<���<K��<2��<���<Z��<w��<���<n��<.��<K��<`   `   ��<A��<���<���<o��<A��<��<���<��<{��<��<���<���<Z��<���<-��<���<Z��<u��<���</��<{��<��<���<`   `   ��<^��<���<���<o��<��<C��<i��<;��<��<���<���<l��<7��<���<p��<��<w��<���<���<n��<2��<p��<R��<`   `   1��<���<��<���<$��< ��<'��<i��<��<n��<F��<���<1��<���<���<���<>��<���</��<n��</��<i��<��< ��<`   `   8��<���<���<5��<���<���<B��<{��<;��<c��<o��<���<��<���<���<��<���<n��<{��<2��<i��<R��<���<���<`   `   ���<���<���<���<���<���<��<p��< ��<.��<���<C��<~��<���<^��<C��<���<.��<��<p��<��<���<���<���<`   `   ���<���<[��<���<���<��<C��<���<T��<���<u��<���<;��<F��<���<u��<���<K��<���<R��< ��<���<���<g��<`   `   ���<���<��<���<N��<Y��<o��<C��<&��<x��<���<���<*��<���<o��<x��<P��<C��<>��<Y��<x��<���<��<���<`   `   ���<[��< ��<���<���<u��<k��<��<��<���<���<-��<!��<���<���<��<���<���<���<���<���<��<b��<���<`   `   ��< ��<v��<K��<]��<��<���<?��<?��<X��<���<a��<���<X��<6��<?��<���<��<Z��<K��<w��< ��<��<C��<`   `   ���<���<K��<-��<���<���<!��<���<��<���<���<���<���<��<���<7��<���<���<G��<\��<���<���<���<���<`   `   N��<���<]��<���<_��<d��<���<e��< ��<���<���<���<:��<e��<\��<d��<���<���<1��<���<h��<���< ��<���<`   `   Y��<u��<��<���<d��<���<5��<���<6��<!��<��<(��<���<K��<���<M��<���<���<���<S��<T��<���<���<g��<`   `   o��<k��<���<!��<���<5��<��<���<n��<F��<~��<���<��<5��<���<!��<���<k��<[��<���<��<V��<���<���<`   `   C��<��<?��<���<e��<���<���<9��<���<���<8��<���<���<N��<���<P��<���<=��<���<���<	��<��<���<t��<`   `   &��<��<?��<��< ��<6��<n��<���<g��<���<Z��<6��<C��<��<��<��<H��<���<���<��<���<��<���<���<`   `   x��<���<X��<���<���<!��<F��<���<���<\��<��<t��<���<j��<���<q��<T��<9��<��<}��<j��<���<@��<p��<`   `   ���<���<���<���<���<��<~��<8��<Z��<��<���<���<���<���<w��<!��<Q��<���<W��<���<���<���<.��<!��<`   `   ���<-��<a��<���<���<(��<���<���<6��<t��<���<r��<!��<���<���<\��<o��<���<��< ��<���<���<b��<���<`   `   *��<!��<���<���<:��<���<��<���<C��<���<���<!��<<��<��<��<���<���<���<?��<���<���<���<��<��<`   `   ���<���<X��<��<e��<K��<5��<N��<��<j��<���<���<��<g��<u��<	��<���<v��<���<���<���<_��<n��<��<`   `   o��<���<6��<���<\��<���<���<���<��<���<w��<���<��<u��<N��<���<:��<!��<��<���<w��<u��<���<���<`   `   x��<��<?��<7��<d��<M��<!��<P��<��<q��<!��<\��<���<	��<���<���<���<���<���<���<���<���<b��<#��<`   `   P��<���<���<���<���<���<���<���<H��<T��<Q��<o��<���<���<:��<���<��<���<6��<���<���<o��<H��<T��<`   `   C��<���<��<���<���<���<k��<=��<���<9��<���<���<���<v��<!��<���<���<��<���<���<���<���<@��<���<`   `   >��<���<Z��<G��<1��<���<[��<���<���<��<W��<��<?��<���<��<���<6��<���<��<��<h��<��<���<���<`   `   Y��<���<K��<\��<���<S��<���<���<��<}��<���< ��<���<���<���<���<���<���<��<���<j��<��<���<���<`   `   x��<���<w��<���<h��<T��<��<	��<���<j��<���<���<���<���<w��<���<���<���<h��<j��<	��<	��<���<T��<`   `   ���<��< ��<���<���<���<V��<��<��<���<���<���<���<_��<u��<���<o��<���<��<��<	��<l��<���<���<`   `   ��<b��<��<���< ��<���<���<���<���<@��<.��<b��<��<n��<���<b��<H��<@��<���<���<���<���<0��<���<`   `   ���<���<C��<���<���<g��<���<t��<���<p��<!��<���<��<��<���<#��<T��<���<���<���<T��<���<���<U��<`   `   +��<���<!��<���<���<���<2��<���<���<:��<���<���<V��<���<��<:��<���<���<���<���<)��<���<��<���<`   `   ���<���<;��<-��<���<���<���<r��<H��<���<���<���<���<���<���<6��<U��<��<���<���<��<R��<���<���<`   `   !��<;��<q��<9��<��<���<���<���<���<���<���<���<���<���<���<���<���<���<��<9��<n��<;��<&��<���<`   `   ���<-��<9��<���<c��<���<��<���<U��<���<.��<3��<���<C��<���<3��<���<F��<���<P��<��<���<���<���<`   `   ���<���<��<c��<��<Z��<b��<1��<��<p��<���<p��<$��<1��<0��<Z��<H��<c��<���<���<��<���<���<���<`   `   ���<���<���<���<Z��<9��<A��<���<���<S��<N��<���<���<\��<P��<>��<���<���<���<y��<��<���<���</��<`   `   2��<���<���<��<b��<A��<���<U��<8��<���<O��<U��<���<A��<h��<��<���<���< ��<���<���<K��<t��<���<`   `   ���<r��<���<���<1��<���<U��<���<���<y��<���<p��<���<��<���<���<U��<���<^��<n��<8��<K��<t��<B��<`   `   ���<H��<���<U��<��<���<8��<���<���<���<"��<���<.��<U��<���<H��<���<���<���<b��<���<b��<��<���<`   `   :��<���<���<���<p��<S��<���<y��<���<���<N��<S��<���<��<���<0��<	��<%��<���<��<��<���<*��<'��<`   `   ���<���<���<.��<���<N��<O��<���<"��<N��<��<.��<���<���<���<h��<���<��<_��<Y��<���<��<���<h��<`   `   ���<���<���<3��<p��<���<U��<p��<���<S��<.��<���<���<���<���<���<��<6��<���<���<#��<,��<���<���<`   `   V��<���<���<���<$��<���<���<���<.��<���<���<���<k��<���<���<���<���<���<x��<���<���<���<���<���<`   `   ���<���<���<C��<1��<\��<A��<��<U��<��<���<���<���<���<���<q��<n��<���<���<���<^��<���<���<���<`   `   ��<���<���<���<0��<P��<h��<���<���<���<���<���<���<���<^��<��<I��<���<��<��<���<���<���<���<`   `   :��<6��<���<3��<Z��<>��<��<���<H��<0��<h��<���<���<q��<��<���<^��<|��<���<��<^��<���<���<m��<`   `   ���<U��<���<���<H��<���<���<U��<���<	��<���<��<���<n��<I��<^��<L��<^��<D��<n��<���<��<���<	��<`   `   ���<��<���<F��<c��<���<���<���<���<%��<��<6��<���<���<���<|��<^��<���<���<���<#��< ��<*��<���<`   `   ���<���<��<���<���<���< ��<^��<���<���<_��<���<x��<���<��<���<D��<���<Q��<���<n��<���<��<^��<`   `   ���<���<9��<P��<���<y��<���<n��<b��<��<Y��<���<���<���<��<��<n��<���<���<^��<��<P��<t��<��<`   `   )��<��<n��<��<��<��<���<8��<���<��<���<#��<���<^��<���<^��<���<#��<n��<��<���<8��<l��<��<`   `   ���<R��<;��<���<���<���<K��<K��<b��<���<��<,��<���<���<���<���<��< ��<���<P��<8��<f��<���<���<`   `   ��<���<&��<���<���<���<t��<t��<��<*��<���<���<���<���<���<���<���<*��<��<t��<l��<���<���<���<`   `   ���<���<���<���<���</��<���<B��<���<'��<h��<���<���<���<���<m��<	��<���<^��<��<��<���<���<���<`   `   >��<���<��<{��<���<���<���<���<��<|��<6��<(��<���<(��<��<|��<C��<���<g��<���<��<{��<���<���<`   `   ���<���<���<��<8��<���<���<���<Q��<���<<��<���<���<C��<���<;��<s��<���<���<��<��<���<���<���<`   `   ��<���<c��<N��<[��<���<p��<���<���<=��<'��<��<)��<=��<���<���<m��<���<a��<N��<Z��<���<��<���<`   `   {��<��<N��<���<���<���<��<���<{��<T��<���<���<L��<e��<���<"��<���<���<��<i��<��<n��<���<���<`   `   ���<8��<[��<���<���<���<���<'��</��<���<��<���<N��<'��<���<���<���<���<&��<8��<���<]��<z��<]��<`   `   ���<���<���<���<���<���<��<���</��<���<���<��<���<*��<���<d��<���<���<���<���<���<I��<L��<���<`   `   ���<���<p��<��<���<��<���<��<���<4��<���<��<���<��<���<��<r��<���<���<���<{��<L��<f��<���<`   `   ���<���<���<���<'��<���<��<s��<9��<#��<l��<#��<���<��<���<���<s��<���<���<J��<T��<e��<M��<���<`   `   ��<Q��<���<{��</��</��<���<9��<`��<9��<���</��<Y��<{��<m��<Q��<:��<��<e��<���<���<���<}��<��<`   `   |��<���<=��<T��<���<���<4��<#��<9��<S��<���<���<L��<W��<���<o��<p��<���<���<���<���<r��<���<���<`   `   6��<<��<'��<���<��<���<���<l��<���<���<*��<���<��<<��<-��<���<���<��<i��<x��<���<��<���<���<`   `   (��<���<��<���<���<��<��<#��</��<���<���< ��<���<��<���<���<���<���<��<���<���<���<���<���<`   `   ���<���<)��<L��<N��<���<���<���<Y��<L��<��<���<��<���<���<���<o �<��<��<��<d �<���<���<���<`   `   (��<C��<=��<e��<'��<*��<��<��<{��<W��<<��<��<���<���<��<��<��<��<�<��<��<���<���<���<`   `   ��<���<���<���<���<���<���<���<m��<���<-��<���<���<��<��<Z�<|�<�<D�<Z�<��<��<x��<���<`   `   |��<;��<���<"��<���<d��<��<���<Q��<o��<���<���<���<��<Z�<��<R�<n�<��<D�<��<���<���<���<`   `   C��<s��<m��<���<���<���<r��<s��<:��<p��<���<���<o �<��<|�<R�<��<R�<w�<��<x �<���<���<p��<`   `   ���<���<���<���<���<���<���<���<��<���<��<���<��<��<�<n�<R�<�<�<��<���<&��<���<���<`   `   g��<���<a��<��<&��<���<���<���<e��<���<i��<��<��<�<D�<��<w�<�<l�<��<s��<���<x��<���<`   `   ���<��<N��<i��<8��<���<���<J��<���<���<x��<���<��<��<Z�<D�<��<��<��<��<���<��<M��<���<`   `   ��<��<Z��<��<���<���<{��<T��<���<���<���<���<d �<��<��<��<x �<���<s��<���< ��<T��<X��<���<`   `   {��<���<���<n��<]��<I��<L��<e��<���<r��<��<���<���<���<��<���<���<&��<���<��<T��<l��<L��<<��<`   `   ���<���<��<���<z��<L��<f��<M��<}��<���<���<���<���<���<x��<���<���<���<x��<M��<X��<L��<���<���<`   `   ���<���<���<���<]��<���<���<���<��<���<���<���<���<���<���<���<p��<���<���<���<���<<��<���<���<`   `   ��<ݼ�<���<���<��<��<���<���<��<���<���<���<O��<���<���<���<8��<���<[��<��<H��<���<m��<ݼ�<`   `   ݼ�<:��<��<d��<���<,��<���<���<c��<���<q��<��<��<z��<��<K��<���<���<E��<v��<T��<��<;��<μ�<`   `   ���<��<5��<-��<��<X��<���<r��<��<��<���<��<���<��<��<r��<���<X��<��<-��<(��<��<���<���<`   `   ���<d��<-��<��<N��<��<���<R��<<��<$��<���<���<��<$��<f��<���<���<+��<*��<I��<T��<���< ��<��<`   `   ��<���<��<N��<���<Y��<*��< ��<���<���<���<���<��< ��<���<Y��<��<N��<���<���<4��<���<���<���<`   `   ��<,��<X��<��<Y��<���<��<��<���<���<���<~��<��<)��<���<6��<���<u��<E��< ��<���<���<���<���<`   `   ���<���<���<���<*��<��<���<���<1��<F��<R��<���<���<��<9��<���<���<���<���<���<���<y��<z��<���<`   `   ���<���<r��<R��< ��<��<���<��<B��<*��<���<���<��<���<f��<���<���<���<e��<���<&��<6��<���<L��<`   `   ��<c��<��<<��<���<���<1��<B��<3��<B��<��<���<��<<��<���<c��</��<���<���<���<���<���<���<���<`   `   ���<���<��<$��<���<���<F��<*��<B��<g��<���<���<��<(��<��<���<L��<7��<"��<|��<l��<	��<7��<g��<`   `   ���<q��<���<���<���<���<R��<���<��<���<���<���<���<q��<���<>��<���<���<���<� �<���<���<o��<>��<`   `   ���<��<��<���<���<~��<���<���<���<���<���<0��<��<y��<q��< �<��<��<l	�<S	�<��<�< �<]��<`   `   O��<��<���<��<��<��<���<��<��<��<���<��<e��<���<��<�	�<��<��<��<��<��<�	�<��<���<`   `   ���<z��<��<$��< ��<)��<��<���<<��<(��<q��<y��<���<�<?�<�<��<f�<�<��<��<+�<�<���<`   `   ���<��<��<f��<���<���<9��<f��<���<��<���<q��<��<?�<�<��<��<:�<��<��</�<?�<��<q��<`   `   ���<K��<r��<���<Y��<6��<���<���<c��<���<>��< �<�	�<�<��<&�<� �<� �<?�<��<��<�	�< �<G��<`   `   8��<���<���<���<��<���<���<���</��<L��<���<��<��<��<��<� �<�!�<� �<��<��<��<��<���<L��<`   `   ���<���<X��<+��<N��<u��<���<���<���<7��<���<��<��<f�<:�<� �<� �<'�<�<�<��<��<7��<���<`   `   [��<E��<��<*��<���<E��<���<e��<���<"��<���<l	�<��<�<��<?�<��<�<v�<l	�<���<"��<���<e��<`   `   ��<v��<-��<I��<���< ��<���<���<���<|��<� �<S	�<��<��<��<��<��<�<l	�<� �<l��<���<���<���<`   `   H��<T��<(��<T��<4��<���<���<&��<���<l��<���<��<��<��</�<��<��<��<���<l��<��<&��<h��<���<`   `   ���<��<��<���<���<���<y��<6��<���<	��<���<�<�	�<+�<?�<�	�<��<��<"��<���<&��<���<���<���<`   `   m��<;��<���< ��<���<���<z��<���<���<7��<o��< �<��<�<��< �<���<7��<���<���<h��<���<���< ��<`   `   ݼ�<μ�<���<��<���<���<���<L��<���<g��<>��<]��<���<���<q��<G��<L��<���<e��<���<���<���< ��<���<`   `   ��<α�<���<��<8��<��<=��<9��<���<���<���<���<&��<���<���<���<���<9��<��<��<g��<��<���<α�<`   `   α�<��<���<���<���<��<G��<���<2��<#��<���<���<���<���<4��<��<���<i��<0��<���<~��<���<��<���<`   `   ���<���<��<���<0��<t��<��<"��<���<K��<��<���<��<K��<���<"��<���<t��<=��<���<��<���<ҵ�<��<`   `   ��<���<���<r��<���<Y��<p��<3��<��<%��<���<���< ��<���<D��<���<A��<]��<���<���<~��<���<_��<`��<`   `   8��<���<0��<���<���<u��<���<s��<��<?��<���<?��<4��<s��<X��<u��<2��<���<���<���<U��<m��<&��<m��<`   `   ��<��<t��<Y��<u��<���<���<K��<S��</��<$��<;��<F��<��<���<R��<A��<���<0��<
��<��<���<���<��<`   `   =��<G��<��<p��<���<���<���<��<��<���<7��<��<���<���<���<p��<���<G��<7��<���<���<Z��<���<���<`   `   9��<���<"��<3��<s��<K��<��<���<���<���<���<1��<F��<Q��<D��<?��<���<)��<���<c��<���<���<b��<���<`   `   ���<2��<���<��<��<S��<��<���<���<���<���<S��<?��<��<���<2��<���<X��<���<���</��<���<��<X��<`   `   ���<#��<K��<%��<?��</��<���<���<���<���<$��<��< ��<h��<4��<���<W��<���<���<*��<��<���<���<o��<`   `   ���<���<��<���<���<$��<7��<���<���<$��<���<���<���<���<���<���<��<h	�<N�<��<q�<h	�<��<���<`   `   ���<���<���<���<?��<;��<��<1��<S��<��<���<��<���<���< �<��<��<��<��<l�<��<��<��<�<`   `   &��<���<��< ��<4��<F��<���<F��<?��< ��<���<���<;��<D�<��<��<��<�#�<A%�<�#�<��<��<��<D�<`   `   ���<���<K��<���<s��<��<���<Q��<��<h��<���<���<D�<��<��<h%�<�*�<�-�<�-�<�*�<[%�<��<��<I�<`   `   ���<4��<���<D��<X��<���<���<D��<���<4��<���< �<��<��<4'�<�.�<�3�<W5�<q3�<�.�<Q'�<��<��< �<`   `   ���<��<"��<���<u��<R��<p��<?��<2��<���<���<��<��<h%�<�.�<5�<9�<9�<+5�<�.�<[%�<��<��<���<`   `   ���<���<���<A��<2��<A��<���<���<���<W��<��<��<��<�*�<�3�<9�<u:�<9�<�3�<�*�<��<��<��<W��<`   `   9��<i��<t��<]��<���<���<G��<)��<X��<���<h	�<��<�#�<�-�<W5�<9�<9�<F5�<�-�<�#�<��<r	�<���<@��<`   `   ��<0��<=��<���<���<0��<7��<���<���<���<N�<��<A%�<�-�<q3�<+5�<�3�<�-�<'%�<��<P�<���<��<���<`   `   ��<���<���<���<���<
��<���<c��<���<*��<��<l�<�#�<�*�<�.�<�.�<�*�<�#�<��<��<��<���<b��<��<`   `   g��<~��<��<~��<U��<��<���<���</��<��<q�<��<��<[%�<Q'�<[%�<��<��<P�<��<T��<���<t��<��<`   `   ��<���<���<���<m��<���<Z��<���<���<���<h	�<��<��<��<��<��<��<r	�<���<���<���<{��<���<J��<`   `   ���<��<ҵ�<_��<&��<���<���<b��<��<���<��<��<��<��<��<��<��<���<��<b��<t��<���<J��<_��<`   `   α�<���<��<`��<m��<��<���<���<X��<o��<���<�<D�<I�< �<���<W��<@��<���<��<��<J��<_��<��<`   `   ���<��<5��<4��<��<���<��<E��<���<��<��<��<	�<��<o�<��<��<E��<���<���<0��<4��<��<��<`   `   ��<O��<���<��<��<���<��<���<���<��<T��<^��<[��<_��<��<���<���<#��<��<��<��<��<M��<ء�<`   `   5��<���<	��<~��<#��<���<���<p��<%��< ��<���<��<���< ��<.��<p��<���<���<1��<~��<���<���<G��<���<`   `   4��<��<~��<���<N��<r��<���<���<5��<`��<��<��<]��<��<���<���<_��</��<���<���<��<%��<F��<H��<`   `   ��<��<#��<N��<���</��<���<���<o��<"��<���<"��<���<���<���</��<��<N��<���<��<��<���<���<���<`   `   ���<���<���<r��</��<���<��<��<[��<"��<��<D��<	��<5��<���<��<_��<���<��<���<��<���<���<!��<`   `   ��<��<���<���<���<��<��<���<Y��<p��<z��<���<���<��<���<���<���<��<��<R��<���<��<���<R��<`   `   E��<���<p��<���<���<��<���<���<���<���<���<���<	��<���<���<���<���<6��<N��<���<��<%��<���<<��<`   `   ���<���<%��<5��<o��<[��<Y��<���<��<���<E��<[��<���<5��<���<���<��<���<#��<���<���<���<6��<���<`   `   ��<��< ��<`��<"��<"��<p��<���<���<���<��<��<]��<:��<��<���<���<��<�<�
�<�
�<��<��<���<`   `   ��<T��<���<��<���<��<z��<���<E��<��<���<��<���<T��<��<�
�<�<��<~�<��<��<��<�<�
�<`   `   ��<^��<��<��<"��<D��<���<���<[��<��<��<��<[��<��<��<>�<c$�<�*�<h-�<V-�<�*�<v$�<;�<��<`   `   	�<[��<���<]��<���<	��<���<	��<���<]��<���<[��<%	�<K�<�"�<�-�<�5�<�;�<=�<�;�<�5�<�-�<�"�<K�<`   `   ��<_��< ��<��<���<5��<��<���<5��<:��<T��<��<K�<�$�<!2�<_=�<�D�<�H�<�H�<�D�<V=�<2�<�$�<N�<`   `   o�<��<.��<���<���<���<���<���<���<��<��<��<�"�<!2�<�?�<J�<�P�<aS�<|P�<J�<@�<!2�<�"�<��<`   `   ��<���<p��<���</��<��<���<���<���<���<�
�<>�<�-�<_=�<J�<�R�<�W�<X�<�R�<J�<V=�<�-�<;�<�
�<`   `   ��<���<���<_��<��<_��<���<���<��<���<�<c$�<�5�<�D�<�P�<�W�<�Y�<�W�<�P�<�D�<�5�<c$�<�<���<`   `   E��<#��<���</��<N��<���<��<6��<���<��<��<�*�<�;�<�H�<aS�<X�<�W�<TS�<�H�<�;�<�*�<��<��<���<`   `   ���<��<1��<���<���<��<��<N��<#��<�<~�<h-�<=�<�H�<|P�<�R�<�P�<�H�<�<�<h-�<~�<�<<��<N��<`   `   ���<��<~��<���<��<���<R��<���<���<�
�<��<V-�<�;�<�D�<J�<J�<�D�<�;�<h-�<��<�
�<���<���<q��<`   `   0��<��<���<��<��<��<���<��<���<�
�<��<�*�<�5�<V=�<@�<V=�<�5�<�*�<~�<�
�<��<��<���<��<`   `   4��<��<���<%��<���<���<��<%��<���<��<��<v$�<�-�<2�<!2�<�-�<c$�<��<�<���<��</��<���<���<`   `   ��<M��<G��<F��<���<���<���<���<6��<��<�<;�<�"�<�$�<�"�<;�<�<��<<��<���<���<���<Է�<F��<`   `   ��<ء�<���<H��<���<!��<R��<<��<���<���<�
�<��<K�<N�<��<�
�<���<���<N��<q��<��<���<F��<ť�<`   `   d��<2��<��<��<���<E��<k��<��<
��<� �<{�<�<S�<�<h�<� �<+��<��<E��<E��<���<��<��<2��<`   `   2��<���<��<<��<���<��<��<u��<���<b��<R��<f�<d�<\��<k��<���<g��<1��<��<k��<5��<.��<���<%��<`   `   ��<��<��<���<��</��<?��<���<���<e��<[��<���<S��<e��<���<���<5��</��<��<���<ܞ�<��<*��<ɐ�<`   `   ��<<��<���<��<U��<^��<��<&��<?��<,��<N��<W��<+��<,��<0��<��<P��<;��<��<��<5��<��<��<��<`   `   ���<���<��<U��<Y��<���<���<:��<���<��<���<��<���<:��<c��<���<���<U��<��<���<���<��<M��<��<`   `   E��<��</��<^��<���<��<���<���<C��<���<���<0��<���<���<$��<���<P��<E��<��<8��<��<���<���<��<`   `   k��<��<?��<��<���<���<��<���<���<*��<���<���<��<���<���<��<8��<��<k��<���<���<X��<���<���<`   `   ��<u��<���<&��<:��<���<���<���<s��<`��<���<���<���< ��<0��<��<g��<��<���<���<���<���<���<���<`   `   
��<���<���<?��<���<C��<���<s��<U��<s��<���<C��<���<?��<���<���<%��<���<��<t��<l��<t��<&��<���<`   `   � �<b��<e��<,��<��<���<*��<`��<s��<C��<���<��<+��<{��<k��<y �<��<R�<��<��<��<��<O�<��<`   `   {�<R��<[��<N��<���<���<���<���<���<���<���<N��<G��<R��<~�<��<$"�<?*�<�.�<%1�</�<?*�<"�<��<`   `   �<f�<���<W��<��<0��<���<���<C��<��<N��<���<d�<�<l"�<;0�<�;�<YC�<�G�<�G�<RC�<�;�<80�<b"�<`   `   S�<d�<S��<+��<���<���<��<���<���<+��<G��<d�<b�<�'�<)9�<�G�<�R�<wZ�<]�<wZ�<�R�<�G�<69�<�'�<`   `   �<\��<e��<,��<:��<���<���< ��<?��<{��<R��<�<�'�<-<�<+N�<�\�<�g�<�l�<�l�<�g�<�\�<!N�<*<�<�'�<`   `   h�<k��<���<0��<c��<$��<���<0��<���<k��<~�<l"�<)9�<+N�<`�<�n�<hw�<�y�<Mw�<�n�<*`�<+N�<+9�<l"�<`   `   � �<���<���<��<���<���<��<��<���<y �<��<;0�<�G�<�\�<�n�<${�<O��<]��<1{�<~n�<�\�<�G�<80�<��<`   `   +��<g��<5��<P��<���<P��<8��<g��<%��<��<$"�<�;�<�R�<�g�<hw�<O��<���<O��<ew�<�g�<�R�<�;�<"�<��<`   `   ��<1��</��<;��<U��<E��<��<��<���<R�<?*�<YC�<wZ�<�l�<�y�<]��<O��<�y�<�l�<xZ�<RC�<I*�<O�<���<`   `   E��<��<��<��<��<��<k��<���<��<��<�.�<�G�<]�<�l�<Mw�<1{�<ew�<�l�<�\�<�G�<�.�<��<,��<���<`   `   E��<k��<���<��<���<8��<���<���<t��<��<%1�<�G�<wZ�<�g�<�n�<~n�<�g�<xZ�<�G�<.1�<��<a��<���<���<`   `   ���<5��<ܞ�<5��<���<��<���<���<l��<��</�<RC�<�R�<�\�<*`�<�\�<�R�<RC�<�.�<��<���<���<���<��<`   `   ��<.��<��<��<��<���<X��<���<t��<��<?*�<�;�<�G�<!N�<+N�<�G�<�;�<I*�<��<a��<���<q��<���<˨�<`   `   ��<���<*��<��<M��<���<���<���<&��<O�<"�<80�<69�<*<�<+9�<80�<"�<O�<,��<���<���<���<j��<��<`   `   2��<%��<ɐ�<��<��<��<���<���<���<��<��<b"�<�'�<�'�<l"�<��<��<���<���<���<��<˨�<��<ސ�<`   `   ah�<�k�<�t�<}��<��<2��<���<L��<���<I	�<��<]"�<�%�<]"�<��<I	�<���<L��<���<2��<��<}��<�t�<�k�<`   `   �k�<q�<@{�<��<��<���<���<d��<���<i��<`�<R�<R�<g�<o��<���<[��<���<���<��<��<O{�<q�<�k�<`   `   �t�<@{�<���<y��<���<���<���<���<���<7��<���<O��<���<7��<���<���<���<���<���<y��<���<@{�<�t�<yr�<`   `   }��<��<y��<	��<��<~��<I��<���<w��<���<��<��<���<j��<���<Z��<v��<���<��<���<��<t��<��<��<`   `   ��<��<���<��<���<\��<l��<���<��<[��<m��<[��<��<���<U��<\��<��<��<���<��<���<~��<��<~��<`   `   2��<���<���<~��<\��<x��<;��<���<���<���<���<{��<���<L��<~��<J��<v��<���<���<)��<C��<���<���<G��<`   `   ���<���<���<I��<l��<;��<���<���<_��<���<s��<���<���<;��<x��<I��<���<���<���<���<v��<���<t��<���<`   `   L��<d��<���<���<���<���<���<���<o��<b��<���<���<���<{��<���<���<[��<C��<���<���<���<���<���<}��<`   `   ���<���<���<w��<��<���<_��<o��<���<o��<U��<���<��<w��<���<���<���<���<L�<��<U�<��<W�<���<`   `   I	�<i��<7��<���<[��<���<���<b��<o��<���<���<J��<���<F��<o��<@	�<��<�<%�<K(�<G(�<%�<�<��<`   `   ��<`�<���<��<m��<���<s��<���<U��<���<���<��<���<`�<��<�(�<f6�<�A�<KH�<�J�<WH�<�A�<`6�<�(�<`   `   ]"�<R�<O��<��<[��<{��<���<���<���<J��<��<^��<R�<T"�<7�<eI�<Y�<�c�<<i�<4i�<�c�<Y�<bI�<�6�<`   `   �%�<R�<���<���<��<���<���<���<��<���<���<R�<�%�<K>�<U�<9i�<�x�<U��<��<U��<�x�<9i�<U�<K>�<`   `   ]"�<g�<7��<j��<���<L��<;��<{��<w��<F��<`�<T"�<K>�<DY�<�q�<:��<���<���<���<���<6��<�q�<BY�<K>�<`   `   ��<o��<���<���<U��<~��<x��<���<���<o��<��<7�<U�<�q�<Ǌ�<���<ȩ�<���<���<���<ъ�<�q�<U�<7�<`   `   I	�<���<���<Z��<\��<J��<I��<���<���<@	�<�(�<eI�<9i�<:��<���<V��<7��<@��<^��<���<6��<9i�<bI�<�(�<`   `   ���<[��<���<v��<��<v��<���<[��<���<��<f6�<Y�<�x�<���<ȩ�<7��<˻�<7��<Ʃ�<���<�x�<Y�<b6�<��<`   `   L��<���<���<���<��<���<���<C��<���<�<�A�<�c�<U��<���<���<@��<7��<���<���<U��<�c�<�A�<�<t��<`   `   ���<���<���<��<���<���<���<���<L�<%�<KH�<<i�<��<���<���<^��<Ʃ�<���<��<<i�<IH�<%�<\�<���<`   `   2��<��<y��<���<��<)��<���<���<��<K(�<�J�<4i�<U��<���<���<���<���<U��<<i�<�J�<G(�<��<���<���<`   `   ��<��<���<��<���<C��<v��<���<U�<G(�<WH�<�c�<�x�<6��<ъ�<6��<�x�<�c�<IH�<G(�<f�<���<g��<C��<`   `   }��<O{�<@{�<t��<~��<���<���<���<��<%�<�A�<Y�<9i�<�q�<�q�<9i�<Y�<�A�<%�<��<���<���<���<l��<`   `   �t�<q�<�t�<��<��<���<t��<���<W�<�<`6�<bI�<U�<BY�<U�<bI�<b6�<�<\�<���<g��<���<��<��<`   `   �k�<�k�<yr�<��<~��<G��<���<}��<���<��<�(�<�6�<K>�<K>�<7�<�(�<��<t��<���<���<C��<l��<��<�r�<`   `   ;�<�?�<L�<�_�<`y�<��< ��<M��<���<��<(�<Y5�<�9�<Y5�<(�<��<���<M��<��<��<hy�<�_�<L�<�?�<`   `   �?�<G�<�T�<ih�<Ȁ�<V��<��<���<��<��<U�<��<��<X�<��<��<���<���<Y��<���<hh�<�T�<G�<�?�<`   `   L�<�T�<pb�<�t�<[��<���<���<���<���<���<a��<���<^��<���<���<���<���<���<`��<�t�<jb�<�T�<L�<I�<`   `   �_�<ih�<�t�<F��<���<��<޹�<���<=��<���<���<���<���<7��<���<��<��<���<I��<�t�<hh�<�_�<4[�<5[�<`   `   `y�<Ȁ�<[��<���<<��<׮�<���<���<)��<R��<b��<R��<.��<���<���<׮�<F��<���<R��<Ȁ�<ey�<�t�<as�<�t�<`   `   ��<V��<���<��<׮�<���<���<���<���<��<{��<���<���<���<���<Ϯ�<��<���<X��<��<���<R��<P��<���<`   `    ��<��<���<޹�<���<���<C��<׽�</��<���<8��<׽�<;��<���<���<޹�<���<��<"��<���<M��<���<M��<���<`   `   M��<���<���<���<���<���<׽�<|��<��<��<y��<߽�<���<���<���<���<���<I��<��<���<���<���<���< ��<`   `   ���<��<���<=��<)��<���</��<��<9��<��<+��<���<0��<=��<���<��<���<�<?	�<,�<�<,�<C	�<�<`   `   ��<��<���<���<R��<��<���<��<��<��<{��<K��<���<���<��<��<�#�<{/�<�8�<�=�<�=�<�8�<y/�<�#�<`   `   (�<U�<a��<���<b��<{��<8��<y��<+��<{��<m��<���<Z��<U�<(�<3>�<�P�<Y_�<�h�<�k�<�h�<Y_�<�P�<3>�<`   `   Y5�<��<���<���<R��<���<׽�<߽�<���<K��<���<���<��<U5�<BQ�<oj�<D�<���<���<���<��<F�<mj�<@Q�<`   `   �9�<��<^��<���<.��<���<;��<���<0��<���<Z��<��<�9�<M[�<�z�<���<���<·�<���<·�<���<���<�z�<M[�<`   `   Y5�<X�<���<7��<���<���<���<���<=��<���<U�<U5�<M[�<��<[��<���<N��<���<���<Q��<���<Y��<��<M[�<`   `   (�<��<���<���<���<���<���<���<���<��<(�<BQ�<�z�<[��<C��<���<���<f��<���<���<F��<[��<�z�<BQ�<`   `   ��<��<���<��<׮�<Ϯ�<޹�<���<��<��<3>�<oj�<���<���<���<���<���<���<���<���<���<���<mj�<7>�<`   `   ���<���<���<��<F��<��<���<���<���<�#�<�P�<D�<���<N��<���<���<��<���<���<N��<���<D�<�P�<�#�<`   `   M��<���<���<���<���<���<��<I��<�<{/�<Y_�<���<·�<���<f��<���<���<d��<���<���<��<\_�<y/�<��<`   `   ��<X��<`��<I��<R��<X��<"��<��<?	�<�8�<�h�<���<���<���<���<���<���<���<���<���<�h�<�8�<F	�<��<`   `   ��<���<�t�<�t�<Ȁ�<��<���<���<,�<�=�<�k�<���<·�<Q��<���<���<N��<���<���<�k�<�=�<&�<���<Ƹ�<`   `   hy�<hh�<jb�<hh�<ey�<���<M��<���<�<�=�<�h�<��<���<���<F��<���<���<��<�h�<�=�<#�<���<G��<���<`   `   �_�<�T�<�T�<�_�<�t�<R��<���<���<,�<�8�<Y_�<F�<���<Y��<[��<���<D�<\_�<�8�<&�<���< ��<P��<�t�<`   `   L�<G�<L�<4[�<as�<P��<M��<���<C	�<y/�<�P�<mj�<�z�<��<�z�<mj�<�P�<y/�<F	�<���<G��<P��<js�<4[�<`   `   �?�<�?�<I�<5[�<�t�<���<���< ��<�<�#�<3>�<@Q�<M[�<M[�<BQ�<7>�<�#�<��<��<Ƹ�<���<�t�<4[�<I�<`   `   E��<X�<x�<.�<�P�<�x�<ڤ�<���<p��<~�<�;�<�M�<)S�<�M�<�;�<~�<k��<���<��<�x�<�P�<.�<|�<X�<`   `   X�<��<j�<�9�<�Z�<�~�<���<7��<���<+	�<f�<�'�<�'�<e�<)	�<���<:��<���<�~�<�Z�< :�<g�<��<Z�<`   `   x�<j�<'2�<{J�<vg�<���<<��<���<���<���<n��<�<n��<���<���<���<=��<���<ug�<{J�<)2�<j�<w�<��<`   `   .�<�9�<{J�<F_�<�v�<��<���<a��<b��<���<���<���<���<e��<^��<���<��<�v�<C_�<xJ�< :�<.�<W(�<W(�<`   `   �P�<�Z�<vg�<�v�<��<`��<Ũ�<���<���<���<@��<���<���<���<˨�<`��<���<�v�<|g�<�Z�<�P�<�J�<~H�<�J�<`   `   �x�<�~�<���<��<`��<i��<P��<1��<��<��<��<��<2��<L��<g��<c��<��<���<�~�<�x�<Eu�<�r�<�r�<Du�<`   `   ڤ�<���<<��<���<Ũ�<P��<���<��<��<���<��<��<���<P��<Ĩ�<���<<��<���<ۤ�<@��<W��<+��<Y��<@��<`   `   ���<7��<���<a��<���<1��<��<��<���<���<��<��<2��<���<^��<���<:��<���<��<~��<x��<v��<~��<���<`   `   p��<���<���<b��<���<��<��<���<���<���<��<��<���<b��<���<���<l��<��<��<��<��<��<��<��<`   `   ~�<+	�<���<���<���<��<���<���<���<���<��<���<���<���<)	�<�<�4�<5F�<�R�<�X�<�X�<�R�<5F�<�4�<`   `   �;�<f�<n��<���<@��<��<��<��<��<��<;��<���<p��<f�<�;�<�X�<�r�<t��<���<���<���<t��<�r�<�X�<`   `   �M�<�'�<�<���<���<��<��<��<��<���<���<�<�'�<�M�<>s�<9��<9��<k��<���<���<m��<6��<8��<@s�<`   `   )S�<�'�<n��<���<���<2��<���<2��<���<���<p��<�'�<&S�<S��<Z��<���<���<���<��<���<���<���<W��<S��<`   `   �M�<e�<���<e��<���<L��<P��<���<b��<���<f�<�M�<S��<���<���<
�<��<H-�<E-�<��<�<���<���<S��<`   `   �;�<)	�<���<^��<˨�<g��<Ĩ�<^��<���<)	�<�;�<>s�<Z��<���<F�<�0�<2G�<�N�<7G�<�0�<B�<���<Z��<>s�<`   `   ~�<���<���<���<`��<c��<���<���<���<�<�X�<9��<���<
�<�0�<\P�<X`�<U`�<YP�<�0�<�<���<8��<�X�<`   `   k��<:��<=��<��<���<��<<��<:��<l��<�4�<�r�<9��<���<��<2G�<X`�<�h�<X`�<2G�<��<���<9��<�r�<�4�<`   `   ���<���<���<�v�<�v�<���<���<���<��<5F�<t��<k��<���<H-�<�N�<U`�<X`�<�N�<E-�<���<m��<s��<5F�<��<`   `   ��<�~�<ug�<C_�<|g�<�~�<ۤ�<��<��<�R�<���<���<��<E-�<7G�<YP�<2G�<E-�<��<���<���<�R�<��<��<`   `   �x�<�Z�<{J�<xJ�<�Z�<�x�<@��<~��<��<�X�<���<���<���<��<�0�<�0�<��<���<���<���<�X�<��<~��<=��<`   `   �P�< :�<(2�< :�<�P�<Eu�<W��<x��<��<�X�<���<m��<���<�<B�<�<���<m��<���<�X�<��<x��<[��<Eu�<`   `   .�<g�<j�<.�<�J�<�r�<+��<v��<��<�R�<t��<6��<���<���<���<���<9��<s��<�R�<��<x��<'��<�r�<�J�<`   `   |�<��<w�<W(�<~H�<�r�<Y��<~��<��<5F�<�r�<8��<W��<���<Z��<8��<�r�<5F�<��<~��<[��<�r�<{H�<W(�<`   `   X�<Z�<��<W(�<�J�<Du�<@��<���<��<�4�<�X�<@s�<S��<S��<>s�<�X�<�4�<��<��<=��<Eu�<�J�<W(�<��<`   `   ���<a��<F��<��<\�<�N�<���<���<���<�.�<�T�<�l�<�t�<�l�<�T�<�.�<���<���<���<�N�<G�<��<R��<a��<`   `   a��<V��<���<���<�%�<�V�<"��<���<���<H�<�*�<�8�<�8�<�*�<A�<���<���<��<�V�<�%�<���<���<W��<h��<`   `   F��<���<���<��<�6�<y`�<8��<G��<��<	��<U�<��<Y�<	��<��<G��<>��<y`�<�6�<��<���<���<=��<���<`   `   ��<���<��<�+�<�J�<(l�<��<2��<?��<���<���<���<���<J��<+��<��<1l�<�J�<�+�<��<���<��<��<��<`   `   \�<�%�<�6�<�J�<Ra�<
y�<���<%��<���<���<���<���<���<%��<���<
y�<:a�<�J�<�6�<�%�<O�<E�<i�<E�<`   `   �N�<�V�<y`�<(l�<
y�<'��<��<���<e��<̥�<ѥ�<p��<���<Ӑ�<!��<y�<1l�<l`�<�V�<�N�<pI�<sF�<tF�<kI�<`   `   ���<"��<8��<��<���<��<:��<���</��<ϗ�<��<���<G��<��<���<��<<��<"��<���<k��<���<j��<���<k��<`   `   ���<���<G��<2��<%��<���<���<���<r��<}��<���<���<���<5��<+��<:��<���<���<���<}��<p��<k��<~��<���<`   `   ���<���<��<?��<���<e��</��<r��<`��<r��<9��<e��<���<?��<.��<���<���<��<��<�$�<�'�<�$�<��<��<`   `   �.�<H�<	��<���<���<̥�<ϗ�<}��<r��<���<ѥ�<���<���<���<A�</�<�J�<�a�<�r�<k{�<o{�<�r�<�a�<�J�<`   `   �T�<�*�<U�<���<���<ѥ�<��<���<9��<ѥ�<���<���<a�<�*�<�T�<[|�<ٞ�<K��<|��<j��<o��<K��<��<[|�<`   `   �l�<�8�<��<���<���<p��<���<���<e��<���<���<��<�8�<�l�<B��<���<���<��<0�<8�<��<���<���<H��<`   `   �t�<�8�<Y�<���<���<���<G��<���<���<���<a�<�8�<�t�<���<���<@�<KD�<�\�<(e�<�\�<PD�<@�<���<���<`   `   �l�<�*�<	��<J��<%��<Ӑ�<��<5��<?��<���<�*�<�l�<���<E��<3�<�e�<S��<���<���<J��<�e�<3�<F��<���<`   `   �T�<A�<��<+��<���<!��<���<+��<.��<A�<�T�<B��<���<3�<�q�<��<���<h��<���<��<�q�<3�<���<B��<`   `   �.�<���<G��<��<
y�<y�<��<:��<���</�<[|�<���<@�<�e�<��<���<��<��<���<��<�e�<?�<���<V|�<`   `   ���<���<>��<1l�<:a�<1l�<<��<���<���<�J�<ٞ�<���<KD�<S��<���<��<0��<��<���<S��<HD�<���<ݞ�<�J�<`   `   ���<��<y`�<�J�<�J�<l`�<"��<���<��<�a�<K��<��<�\�<���<h��<��<��<n��<���<�\�<��<F��<�a�<��<`   `   ���<�V�<�6�<�+�<�6�<�V�<���<���<��<�r�<|��<0�<(e�<���<���<���<���<���<1e�<0�<}��<�r�<��<���<`   `   �N�<�%�<��<��<�%�<�N�<k��<}��<�$�<k{�<j��<9�<�\�<J��<��<��<S��<�\�<0�<e��<o{�<�$�<~��<\��<`   `   G�<���<���<���<O�<pI�<���<p��<�'�<o{�<o��<��<PD�<�e�<�q�<�e�<HD�<��<}��<o{�<�'�<p��<É�<pI�<`   `   ��<���<���<��<E�<sF�<j��<k��<�$�<�r�<K��<���<@�<3�<3�<?�<���<F��<�r�<�$�<p��<[��<tF�<U�<`   `   R��<W��<=��<��<i�<tF�<���<~��<��<�a�<��<���<���<F��<���<���<ݞ�<�a�<��<~��<É�<tF�<X�<��<`   `   a��<h��<���<��<E�<kI�<k��<���<��<�J�<[|�<H��<���<���<B��<V|�<�J�<��<���<\��<pI�<U�<��<���<`   `   �7�<=B�<}_�<��<���<��<�b�<Բ�<c��<�@�<�s�<7��<���<7��<�s�<�@�<A��<Բ�<�b�<��<���<��<�_�<=B�<`   `   =B�<�R�<�s�<��<a��<>�<�b�<���<���<��<�;�<�N�<�N�<�;�<��<���<���<�b�<0�<{��<���<qs�<�R�<KB�<`   `   }_�<�s�<��<_��<z��<�+�<�d�<���<���<q��<��<��<��<q��<���<���<�d�<�+�<n��<_��< ��<�s�<m_�<{X�<`   `   ��<��<_��<���<��<�;�<&g�<)��<1��<���< ��<���<���<D��<��<g�<�;�<��<���<I��<���< ��<3��<1��<`   `   ���<a��<z��<��<M-�<�L�<rj�<ф�<��<6��<���<6��<ܘ�<ф�<�j�<�L�<#-�<��<���<a��<���<��<��<��<`   `   ��<>�<�+�<�;�<�L�<a^�<�n�<0|�<?��<I��<R��<R��<2|�<�n�<V^�<�L�<�;�<�+�<0�<��<��<��<��<��<`   `   �b�<�b�<�d�<&g�<rj�<�n�<Kr�<>u�<�w�<�w�<�w�<>u�<cr�<�n�<bj�<&g�<�d�<�b�<�b�<b�<=b�<Nb�<Bb�<b�<`   `   Բ�<���<���<)��<ф�<0|�<>u�<|q�<o�<o�<�q�<$u�<2|�<��<��<y��<���<��<Ӽ�<K��<0��<)��<M��<��<`   `   c��<���<���<1��<��<?��<�w�<o�<�k�<o�<�w�<?��<Ԙ�<1��<��<���<G��<��<�'�<�3�<J7�<�3�<�'�<��<`   `   �@�<��<q��<���<6��<I��<�w�<o�<o�<�w�<R��<P��<���<[��<��<�@�< f�<���<���<;��<B��<���<���<f�<`   `   �s�<�;�<��< ��<���<R��<�w�<�q�<�w�<R��<���< ��<��<�;�<�s�<#��<���<]��<��<��<��<]��<��<#��<`   `   7��<�N�<��<���<6��<R��<>u�<$u�<?��<P��< ��<��<�N�<D��<���<O�<�K�<�p�<���<���<q�<zK�<R�<���<`   `   ���<�N�<��<���<ܘ�<2|�<cr�<2|�<Ԙ�<���<��<�N�<���<���<�?�<3��<s��<!��<p��<!��<z��<3��<w?�<���<`   `   7��<�;�<q��<D��<ф�<�n�<�n�<��<1��<[��<�;�<D��<���<xM�<¡�<��<��<<3�<.3�<��<$��<͡�<zM�<���<`   `   �s�<��<���<��<�j�<V^�<bj�<��<��<��<�s�<���<�?�<¡�<���<|9�<c�<�q�<�c�<|9�<���<¡�<�?�<���<`   `   �@�<���<���<g�<�L�<�L�<&g�<y��<���<�@�<#��<O�<3��<��<|9�<gt�<���<���<Yt�<�9�<$��<2��<R�<��<`   `   A��<���<�d�<�;�<#-�<�;�<�d�<���<G��< f�<���<�K�<s��<��<c�<���<c��<���<�c�<��<m��<�K�<��< f�<`   `   Բ�<�b�<�+�<��<��<�+�<�b�<��<��<���<]��<�p�<!��<<3�<�q�<���<���< r�<.3�<��<q�<T��<���<��<`   `   �b�<0�<n��<���<���<0�<�b�<Ӽ�<�'�<���<��<���<p��<.3�<�c�<Yt�<�c�<.3�<���<���<��<���<�'�<Ӽ�<`   `   ��<{��<_��<I��<a��<��<b�<K��<�3�<;��<��<���<!��<��<|9�<�9�<��<��<���<��<B��<�3�<M��<�a�<`   `   ���<���< ��<���<���<��<=b�<0��<J7�<B��<��<q�<z��<$��<���<$��<m��<q�<��<B��</7�<0��<Tb�<��<`   `   ��<qs�<�s�< ��<��<��<Nb�<)��<�3�<���<]��<zK�<3��<͡�<¡�<2��<�K�<T��<���<�3�<0��<5b�<��<���<`   `   �_�<�R�<m_�<3��<��<��<Bb�<M��<�'�<���<��<R�<w?�<zM�<�?�<R�<��<���<�'�<M��<Tb�<��<Ѽ�<3��<`   `   =B�<KB�<{X�<1��<��<��<b�<��<��<f�<#��<���<���<���<���<��< f�<��<Ӽ�<�a�<��<���<3��<dX�<`   `   0��<C��<B��<��<�a�<���<s+�</��<y��<DV�<���<���<��<���<қ�<DV�<J��</��<�+�<���<�a�<��<]��<C��<`   `   C��<��<��<H,�<5y�<���<�,�<��<���<b�<�P�<j�<j�<�P�<S�<��<4��<�,�<���<Yy�<S,�<���<��<U��<`   `   B��<��<R�<cS�<]��<���<�/�<�w�<��<w��<0�<��<9�<w��<��<�w�<�/�<���<L��<cS�<e�<��<-��<���<`   `   ��<H,�<cS�<q��<��<V��<�2�<�h�<��<��<F��<:��<��<��<�h�<}2�<k��</��<]��<ES�<S,�<�<@�<=�<`   `   �a�<5y�<]��<��<���<�<	8�<�\�<�w�<��<P��<��<w�<�\�<:8�<�<t��<��<���<5y�<�a�<�S�<�N�<�S�<`   `   ���<���<���<V��<�<2(�<�=�<�Q�<_�<�f�<�f�<_�<�Q�<�=�<#(�<:�<k��<���<���<���<���<���<���<���<`   `   s+�<�,�<�/�<�2�<	8�<�=�<D�<|I�<{M�<�N�<UM�<|I�<5D�<�=�<�7�<�2�<�/�<�,�<u+�<v+�<�+�<f+�<�+�<v+�<`   `   /��<��<�w�<�h�<�\�<�Q�<|I�<iE�<�B�<�B�<vE�<YI�<�Q�<�\�<�h�<�w�<4��<A��<k��<���<���<���<���<��<`   `   y��<���<��<��<�w�<_�<{M�<�B�<�=�<�B�<�M�<_�<uw�<��<D��<���<R��<(�<;4�<�C�<bI�<�C�<$4�<(�<`   `   DV�<b�<w��<��<��<�f�<�N�<�B�<�B�<eN�<�f�<;��<��<Y��<S�<VV�<ӈ�<޳�<P��<W��<b��<d��<��<���<`   `   ���<�P�<0�<F��<P��<�f�<UM�<vE�<�M�<�f�< ��<F��<K�<�P�<���<X��<�"�<*T�<�s�<�~�<�s�<*T�<�"�<X��<`   `   ���<j�<��<:��<��<_�<|I�<YI�<_�<;��<F��<p�<j�<���<O$�<Jy�<��<2��<�<�<=��<Կ�<Ly�<^$�<`   `   ��<j�<9�<��<w�<�Q�<5D�<�Q�<uw�<��<K�<j�<���<�E�<k��<��<�V�<K��<֔�<K��<�V�<��<Y��<�E�<`   `   ���<�P�<w��<��<�\�<�=�<�=�<�\�<��<Y��<�P�<���<�E�<���<�5�<l��<d��<f��<S��<O��<w��<�5�<���<�E�<`   `   қ�<S�<��<�h�<:8�<#(�<�7�<�h�<D��<S�<���<O$�<k��<�5�<��<'�<-A�</U�<VA�<'�<ת�<�5�<k��<O$�<`   `   DV�<��<�w�<}2�<�<:�<�2�<�w�<���<VV�<X��<Jy�<��<l��<'�<rX�<���<k��<^X�<6�<w��<��<Ly�<L��<`   `   J��<4��<�/�<k��<t��<k��<�/�<4��<R��<ӈ�<�"�<��<�V�<d��<-A�<���<���<���<2A�<d��<�V�<��<�"�<ӈ�<`   `   /��<�,�<���</��<��<���<�,�<A��<(�<޳�<*T�<2��<K��<f��</U�<k��<���<>U�<S��<H��<=��<T�<��<B�<`   `   �+�<���<L��<]��<���<���<u+�<k��<;4�<P��<�s�<�<֔�<S��<VA�<^X�<2A�<S��<��<�<�s�<P��<4�<k��<`   `   ���<Yy�<cS�<ES�<5y�<���<v+�<���<�C�<W��<�~�<�<K��<O��<'�<6�<d��<H��<�<�~�<b��<�C�<���<S+�<`   `   �a�<S,�<e�<S,�<�a�<���<�+�<���<bI�<b��<�s�<=��<�V�<w��<ת�<w��<�V�<=��<�s�<b��<>I�<���< ,�<���<`   `   ��<���<��<�<�S�<���<f+�<���<�C�<d��<*T�<Կ�<��<�5�<�5�<��<��<T�<P��<�C�<���<C+�<���<�S�<`   `   ]��<��<-��<@�<�N�<���<�+�<���<$4�<��<�"�<Ly�<Y��<���<k��<Ly�<�"�<��<4�<���< ,�<���<[N�<@�<`   `   C��<U��<���<=�<�S�<���<v+�<��<(�<���<X��<^$�<�E�<�E�<O$�<L��<ӈ�<B�<k��<S+�<���<�S�<@�<o��<`   `   ���<���<6�<�g�<���<�R�<���<�n�<���<(p�<,��<	�<�<	�<M��<(p�<|��<�n�<-��<�R�<}��<�g�<X�<���<`   `   ���<D�<�:�<���<W��<�f�<���<AZ�<.��<�&�<i�<���<��<i�<�&�<M��<\Z�<���<xf�<���<���<x:�<G�<���<`   `   6�<�:�<ft�<p��<U�<�~�<d��<�F�<���<x��<@	�<��<I	�<x��<���<�F�<r��<�~�<C�<p��<{t�<�:�< �<�
�<`   `   �g�<���<p��<D�<�L�<���<}��<4�<jp�<]��<���<s��<a��<�p�<�3�<T��<��<
M�<+�<L��<���<�g�<�U�<�U�<`   `   ���<W��<U�<�L�<^��<=��<~��<�#�<4J�<�b�<�j�<�b�<J�<�#�<���<=��<��<�L�<��<W��<���<x��< ��<x��<`   `   �R�<�f�<�~�<���<=��<���<���<!�<�+�<W5�<e5�<�+�<&�<���<���<h��<��<�~�<xf�<�R�<�E�<&?�<(?�<�E�<`   `   ���<���<d��<}��<~��<���<�<b�<��<�<��<b�<*�<���<g��<}��<m��<���<���<?��<���<5��<���<?��<`   `   �n�<AZ�<�F�<4�<�#�<!�<b�<��<!�<?�<��<9�<&�<�#�<�3�<`F�<\Z�<�n�<���<ۍ�<��<Ԕ�<ލ�<Հ�<`   `   ���<.��<���<jp�<4J�<�+�<��<!�<��<!�<��<�+�<J�<jp�<��<.��<���< !�<PA�<�V�<�^�<�V�<4A�< !�<`   `   (p�<�&�<x��<]��<�b�<W5�<�<?�<!�<��<e5�<*c�<a��<T��<�&�<<p�<��<���<E�<�-�<�-�<^�<���<س�<`   `   ,��<i�<@	�<���<�j�<e5�<��<��<��<e5�<�j�<���<_	�<i�<+��<�.�<ڄ�<_��<���<c�<r��<_��<��<�.�<`   `   	�<���<��<s��<�b�<�+�<b�<9�<�+�<*c�<���<��<��<-	�<��<?��<p[�<���<{��<���<���<U[�<B��<%��<`   `   �<��<I	�<a��<J�<&�<*�<&�<J�<a��<_	�<��<��<j��<E�<,��<�)�<�i�<��<�i�<�)�<,��<E�<j��<`   `   	�<i�<x��<�p�<�#�<���<���<�#�<jp�<T��<i�<-	�<j��<�^�<���<o��<S��<[�<B�<8��<~��<���<�^�<e��<`   `   M��<�&�<���<�3�<���<���<g��<�3�<��<�&�<+��<��<E�<���<��<�<�m�<(��<�m�<�<]��<���<E�<��<`   `   (p�<M��<�F�<T��<=��<h��<}��<`F�<.��<<p�<�.�<?��<,��<o��<�<Q��<���<w��<8��<$�<~��<(��<B��<.�<`   `   |��<\Z�<r��<��<��<��<m��<\Z�<���<��<ڄ�<p[�<�)�<S��<�m�<���<L��<���<�m�<S��<�)�<p[�<��<��<`   `   �n�<���<�~�<
M�<�L�<�~�<���<�n�< !�<���<_��<���<�i�<\�<(��<w��<���<<��<B�<�i�<���<R��<���<!�<`   `   -��<xf�<C�<+�<��<xf�<���<���<PA�<E�<���<{��<��<B�<�m�<8��<�m�<B�<��<{��<���<E�</A�<���<`   `   �R�<���<o��<L��<W��<�R�<?��<ۍ�<�V�<�-�<c�<���<�i�<8��<�<$�<S��<�i�<{��<U�<�-�<�V�<ލ�<��<`   `   }��<���<{t�<���<���<�E�<���<��<�^�<�-�<r��<���<�)�<~��<]��<~��<�)�<���<���<�-�<n^�<��<���<�E�<`   `   �g�<x:�<�:�<�g�<x��<&?�<5��<Ԕ�<�V�<^�<_��<U[�<,��<���<���<(��<p[�<R��<E�<�V�<��<��<(?�<���<`   `   X�<G�< �<�U�< ��<(?�<���<ލ�<4A�<���<��<B��<E�<�^�<E�<B��<��<���</A�<ލ�<���<(?�<ӹ�<�U�<`   `   ���<���<�
�<�U�<x��<�E�<?��<Հ�< !�<س�<�.�<%��<j��<e��<��<.�<��<!�<���<��<�E�<���<�U�<�
�<`   `   ���<���<��<K��<I�<[��<t�<�4�<��<R��<q�<`]�<y�<`]�<��<R��<���<�4�<�t�<[��<�<K��<��<���<`   `   ���<���<bJ�<��<!;�<z��<+x�<�<O��<a-�<j��<���<���<]��<I-�<o��<;�<�w�<[��<P;�<%��<;J�<���<���<`   `   ��<bJ�<_��<���<\q�<��<:�<� �<�s�<T��<�<��<�<T��<�s�<� �<F�<��<Kq�<���<s��<bJ�<{�<��<`   `   K��<��<���<�P�<��<��<���<��<%<�<�v�<s��<e��<�v�<F<�<��<���<��<��<�P�<���<%��<`��<�l�<�l�<`   `   I�< ;�<\q�<��<���<4K�<2��<X��<��<�-�<G8�<�-�<f�<X��<w��<4K�<q��<��<�q�< ;�<!�<*��<���<*��<`   `   [��<z��<��<��<4K�<�y�<���<"��< ��<"��<0��<A��<)��<m��<�y�<cK�<��<���<[��<q��<)��<%��<&��<��<`   `   t�<+x�<:�<���<2��<���<��<Y��<���<���<���<Y��<��<���<��<���<@�<+x�<�t�<�r�<Cs�<�r�<Ts�<�r�<`   `   �4�<�<� �<��<X��<"��<Y��<V��<���<���<d��<,��<)��<���<��<� �<;�<�4�<�K�<�\�<Af�</f�<�\�<�K�<`   `   ��<N��<�s�<%<�<��< ��<���<���<ô�<���<��< ��<W�<%<�<4t�<N��<���<�"�<�N�<3k�<�t�<3k�<�N�<�"�<`   `   R��<a-�<T��<�v�<�-�<"��<���<���<���<���<0��<�-�<�v�<-��<I-�<h��<���<�6�<�o�<���<Ҍ�<�o�<�6�<���<`   `   q�<j��<�<s��<G8�<0��<���<d��<��<0��<
8�<s��<%�<j��<t�<<��<�<`�<��<���<O��<`�<"�<<��<`   `   `]�<���<��<e��<�-�<A��<Y��<,��< ��<�-�<s��<[�<���<v]�<��<ʤ�<�)�<h��<���<ý�<{��<�)�<ˤ�<��<`   `   y�<���<�<�v�<f�<)��<��<)��<W�<�v�<%�<���<�x�<9E�<M�<��<�F�<���<A��<���<�F�<��<4�<9E�<`   `   `]�<]��<T��<F<�<X��<m��<���<���<%<�<-��<j��<v]�<9E�<�.�<��<���<�B�<���<���<�B�<���<��<�.�<2E�<`   `   ��<I-�<�s�<��<w��<�y�<��<��<4t�<I-�<t�<��<M�<��<���<̘�<�	�<�0�<�	�<̘�<���<��<S�<��<`   `   R��<o��<� �<���<4K�<cK�<���<� �<N��<h��<<��<ʤ�<��<���<̘�<�6�<��<��<�6�<��<���<x��<ˤ�</��<`   `   ���<;�<F�<��<q��<��<@�<;�<���<���<�<�)�<�F�<�B�<�	�<��<1��<��<�	�<�B�<�F�<�)�<�<���<`   `   �4�<�w�<��<��<��<���<+x�<�4�<�"�<�6�<`�<h��<���<���<�0�<��<��<�0�<���<���<{��<`�<�6�<#�<`   `   �t�<[��<Kq�<�P�<�q�<[��<�t�<�K�<�N�<�o�<��<���<A��<���<�	�<�6�<�	�<���<g��<���<{��<�o�<�N�<�K�<`   `   [��<P;�<���<���< ;�<q��<�r�<�\�<3k�<���<���<ý�<���<�B�<̘�<��<�B�<���<���<���<Ҍ�<Sk�<�\�<�r�<`   `   �<%��<s��<%��<!�<)��<Cs�<Af�<�t�<Ҍ�<O��<{��<�F�<���<���<���<�F�<{��<{��<Ҍ�<rt�<Af�<os�<)��<`   `   K��<;J�<bJ�<`��<*��<%��<�r�</f�<3k�<�o�<`�<�)�<��<��<��<x��<�)�<`�<�o�<Sk�<Af�<�r�<&��<Y��<`   `   ��<���<{�<�l�<���<&��<Ts�<�\�<�N�<�6�<"�<ˤ�<4�<�.�<S�<ˤ�<�<�6�<�N�<�\�<os�<&��<���<�l�<`   `   ���<���<��<�l�<*��<��<�r�<�K�<�"�<���<=��<��<9E�<2E�<��</��<���<#�<�K�<�r�<)��<Y��<�l�<��<`   `   n\�<Ky�<���<�V�<��<���<��<���<d��<���<�Y�<9��<���<9��<Z�<���<��<���<S��<���<J�<�V�<��<Ky�<`   `   Ky�<$��<W
�<��<�D�<��<���<��<;��<�.�<���<��< ��<��<�.�<\��<��<i��<g�<�D�<"��<0
�<#��<`y�<`   `   ���<W
�<�l�<��<���<�<�<���<���<�9�<���<, �<��<. �<���<�9�<���<���<�<�<���<��<�l�<W
�<���<]��<`   `   �V�<��<��<c�<���<�t�<�<���<E��<C�<1m�<%m�< C�<f��<���<��<�t�<���<�b�<���<"��<�V�<�6�<�6�<`   `   ��<�D�<���<���<&K�<d��<��<�r�<޸�<���<���<���<���<�r�<�<d��<�J�<���<��<�D�<e�<Y��<���<Y��<`   `   ���<��<�<�<�t�<d��<��<60�<�d�<9��<S��<`��<Z��<�d�<	0�<���<���<�t�<�<�<g�<���<���<���<���<}��<`   `   ��<���<���<�<��<60�<_H�<�\�<k�<�n�<�j�<�\�<�H�<60�<��<�<���<���<��<d��<���<p��<���<d��<`   `   ���<��<���<���<�r�<�d�<�\�<�Y�<_W�<W�<�Y�<�\�<�d�<s�<���<w��<��<���<{��<H�<��<��<G�<���<`   `   d��<;��<�9�<E��<޸�<9��<k�<_W�<wP�<_W�<$k�<9��<���<E��<�9�<;��<*��<:�<9W�<~�<P��<~�<W�<:�<`   `   ���<�.�<���<C�<���<S��<�n�<W�<_W�<un�<`��<���< C�<{��<�.�<ͮ�<M)�<��<��<��<��<3��<��<()�<`   `   �Y�<���<, �<1m�<���<`��<�j�<�Y�<$k�<`��<H��<1m�<I �<���<�Y�<
�<���<�!�<�s�<��<�s�<�!�<���<
�<`   `   9��<��<��<%m�<���<Z��<�\�<�\�<9��<���<1m�<{�< ��<N��<­�<��<�6�<P��<,�<O�<f��<�6�<��<ݭ�<`   `   ���< ��<. �< C�<���<�d�<�H�<�d�<���< C�<I �< ��<���<���<��<���<��<j<�<g�<j<�<��<���<j�<���<`   `   9��<��<���<f��<�r�<	0�<60�<s�<E��<{��<���<N��<���<1=�<=i�<�f�<��<V��<4��<��<g�<Xi�</=�<���<`   `   Z�<�.�<�9�<���<�<���<��<���<�9�<�.�<�Y�<­�<��<=i�<A��<��<g5�<�k�<�5�<��<��<=i�<��<­�<`   `   ���<\��<���<��<d��<���<�<w��<;��<ͮ�<
�<��<���<�f�<��<�t�<���<���<ot�<9��<g�<���<��<
�<`   `   ��<��<���<�t�<�J�<�t�<���<��<*��<M)�<���<�6�<��<��<g5�<���<�%�<���<n5�<��<��<�6�<���<M)�<`   `   ���<i��<�<�<���<���<�<�<���<���<:�<��<�!�<P��<j<�<V��<�k�<���<���<l�<4��<`<�<f��<�!�<��<Z�<`   `   S��<g�<���<�b�<��<g�<��<{��<9W�<��<�s�<,�<g�<4��<�5�<ot�<n5�<4��<4g�<,�<�s�<��<W�<{��<`   `   ���<�D�<��<���<�D�<���<d��<H�<~�<��<��<O�<j<�<��<��<9��<��<`<�<,�< ��<��<;~�<G�<6��<`   `   J�<"��<�l�<"��<e�<���<���<��<P��<��<�s�<f��<��<g�<��<g�<��<f��<�s�<��<��<��<���<���<`   `   �V�<0
�<W
�<�V�<Y��<���<p��<��<~�<3��<�!�<�6�<���<Xi�<=i�<���<�6�<�!�<��<;~�<��<B��<���<���<`   `   ��<#��<���<�6�<���<���<���<G�<W�<��<���<��<j�</=�<��<��<���<��<W�<G�<���<���<���<�6�<`   `   Ky�<`y�<]��<�6�<Y��<}��<d��<���<:�<()�<
�<ݭ�<���<���<­�<
�<M)�<Z�<{��<6��<���<���<�6�<6��<`   `   ���<���<��<���<���<��<��<�]�<x��<���<T��<mF�<�y�<mF�<|��<���<3��<�]�<�<��<J��<���<��<���<`   `   ���<~��<�b�<��<���<� �<��<�;�<3B�<#�<���<K�<X�<���<�"�<PB�<<�<��<� �<!��<��<�b�<z��<���<`   `   ��<�b�<l��<��<�[�<SA�<�1�<��<>��<���<���<�<���<���<?��<��<�1�<SA�<�[�<��<w��<�b�<��<���<`   `   ���<��<��<�$�<��<���<�L�<V��<A��< ��<�2�<�2�<-��<^��<7��<�L�<��<I��<�$�<͌�<��<���<ՙ�<ٙ�<`   `   ���<���<�[�<��<Y�<$��<o�<4��<sI�<���<˜�<���<II�<4��<Zo�<$��<�X�<��<�[�<���<e��<���<�t�<���<`   `   ��<� �<SA�<���<$��<�@�<u��<8��<��<�1�<�1�<��<E��<J��<w@�<Q��<��</A�<� �<��<���<���<���<���<`   `   ��<��<�1�<�L�<o�<u��<���<t��<��<��<���<t��<���<u��<o�<�L�<�1�<��<��<C�<��<�<�<C�<`   `   �]�<�;�<��<V��<4��<8��<t��<S��<b��<��<\��<I��<E��<a��<7��<��<<�<�]�<d��<���<��<���<���<���<`   `   x��<3B�<>��<A��<sI�<��<��<b��<	��<b��<@��<��<:I�<A��<���<3B�<>��<i�<UP�<��<���<��<4P�<i�<`   `   ���<#�<���< ��<���<�1�<��<��<b��<���<�1�<ч�<-��<b��<�"�<���<�l�<c��<�]�<���<ѓ�<^�<_��<gl�<`   `   T��<���<���<�2�<˜�<�1�<���<\��<@��<�1�<���<�2�<���<���<a��<��<Kq�<��<n��<��<0��<��<wq�<��<`   `   mF�<K�<�<�2�<���<��<t��<I��<��<ч�<�2�<��<X�<F�<Zy�<v��<��<�F�< ��<%��<G�<ɒ�<r��<yy�<`   `   �y�<X�<���<-��<II�<E��<���<E��<:I�<-��<���<X�<ry�<Z��<�Z�<f��<ը�<�O�<Q��<�O�<��<f��<�Z�<Z��<`   `   mF�<���<���<^��<4��<J��<u��<a��<A��<b��<���<F�<Z��<P��<W3�<���<���<	�<��<���<��<v3�<L��<M��<`   `   |��<�"�<?��<7��<Zo�<w@�<o�<7��<���<�"�<a��<Zy�<�Z�<W3�<���<�'�<���<�H�<8��<�'�<g��<W3�<�Z�<Zy�<`   `   ���<PB�<��<�L�<$��<Q��<�L�<��<3B�<���<��<v��<f��<���<�'�<+S�<���<h��<S�<�'�<��<Z��<r��<v��<`   `   3��<<�<�1�<��<�X�<��<�1�<<�<>��<�l�<Kq�<��<ը�<���<���<���<AE�<���<���<���<ɨ�<��<Yq�<�l�<`   `   �]�<��<SA�<I��<��</A�<��<�]�<i�<d��<��<�F�<�O�<	�<�H�<h��<���<�H�<��<�O�<G�<��<_��<��<`   `   �<� �<�[�<�$�<�[�<� �<��<d��<UP�<�]�<n��< ��<Q��<��<8��<S�<���<��<���< ��<^��<�]�<;P�<d��<`   `   ��<!��<��<͌�<���<��<C�<���<��<���<��<%��<�O�<���<�'�<�'�<���<�O�< ��<��<ѓ�<-��<���<�<`   `   J��<��<w��<��<e��<���<��<��<���<ѓ�<0��<G�<��<��<h��<��<ɨ�<G�<^��<ѓ�<b��<��<�<���<`   `   ���<�b�<�b�<���<���<���<�<���<��<^�<��<ɒ�<f��<v3�<W3�<Z��<��<��<�]�<-��<��<��<���<���<`   `   ��<z��<��<ՙ�<�t�<���<�<���<4P�<_��<wq�<r��<�Z�<L��<�Z�<r��<Yq�<_��<<P�<���<�<���<�t�<ՙ�<`   `   ���<���<���<ٙ�<���<���<C�<���<i�<gl�<��<yy�<Z��<M��<Zy�<v��<�l�<��<d��<�<���<���<ՙ�<���<`   `   :�<�K�<���<خ�<���<}G�<���</��<�P�<���<���<��<��<��< �<���<ZP�</��<��<}G�<@��<خ�<���<�K�<`   `   �K�<���<�5�<��<�=�<���<��<)y�<���<`�<���<�I�<J�<���<@�<���<Ry�<n�<Ӎ�<
>�<��<�5�<���<	L�<`   `   ���<�5�<1��<@��<���<W��<`$�<�U�<ge�<�<�<��<���<��<�<�<oe�<�U�<\$�<W��<���<@��<5��<�5�<���<��<`   `   خ�<��<@��<�|�<�d�<n\�<�R�<�<�<d�<א�<C��<=��<��<|�<�<�<�R�<�\�<�d�<�|�<!��<��<��<�w�<�w�<`   `   ���<�=�<���<�d�<O�<���<��<&5�<��<��<4#�<��<ŵ�<&5�<9��<���< �<�d�<��<�=�<Z��<���<e��<���<`   `   }G�<���<W��<n\�<���<U�<���<�3�<��<��<��<��<�3�<���<�T�<���<�\�<9��<Ӎ�<�G�<��<�<�<��<`   `   ���<��<`$�<�R�<��<���<��<�9�<7[�<�f�<[�<�9�<��<���<��<�R�<V$�<��<���<���<���<���<���<���<`   `   /��<)y�<�U�<�<�<&5�<�3�<�9�<�A�<G�< G�<�A�<�9�<�3�<M5�<�<�<aU�<Ry�<<��<q��<y��<��<���<r��<���<`   `   �P�<���<ge�<d�<��<��<7[�<G�<�?�<G�<V[�<��<���<d�<�e�<���<eP�<���<��<�W�<�l�<�W�<��<���<`   `   ���<`�<�<�<א�<��<��<�f�< G�<G�<yf�<��<�<��<v<�<@�<���<���<�@�<���<M �<g �<��<�@�<̕�<`   `   ���<���<��<C��<4#�<��<[�<�A�<V[�<��<#�<C��<,��<���<  �<1$�<�+�<���<6��<���<���<���<�+�<1$�<`   `   ��<�I�<���<=��<��<��<�9�<�9�<��<�<C��<���<J�<��<CD�<��<5��<���<g;�<�;�<���<��<��<cD�<`   `   ��<J�<��<��<ŵ�<�3�<��<�3�<���<��<+��<J�<��<���<���<�E�<���<6^�<g��<6^�<���<�E�<ߨ�<���<`   `   ��<���<�<�<|�<&5�<���<���<M5�<d�<v<�<���<��<���<���<��<[��<p��<���<x��<H��<v��<3��<���<{��<`   `    �<@�<oe�<�<�<9��<�T�<��<�<�<�e�<@�<  �<CD�<���<��<,�<��<��<�+�<i��<��<��<��<��<CD�<`   `   ���<���<�U�<�R�<���<���<�R�<aU�<���<���<1$�<��<�E�<[��<��<�:�<��<f�<�:�<4��<v��<E�<��<+$�<`   `   ZP�<Ry�<\$�<�\�< �<�\�<V$�<Ry�<eP�<���<�+�<6��<���<p��<��<��<Yo�<��< ��<p��<���<6��<�+�<���<`   `   /��<n�<W��<�d�<�d�<9��<��<<��<���<�@�<���<���<6^�<���<�+�<f�<��<�+�<x��<&^�<���<���<�@�<���<`   `   ��<Ӎ�<���<�|�<��<Ӎ�<���<q��<��<���<6��<g;�<g��<x��<i��<�:�< ��<x��<���<g;�<!��<���<��<q��<`   `   }G�<
>�<@��<!��<�=�<�G�<���<y��<�W�<M �<���<�;�<6^�<H��<��<4��<p��<&^�<g;�<���<g �<X�<r��<���<`   `   @��<��<5��<��<Z��<��<���<��<�l�<g �<���<���<���<v��<��<v��<���<���<!��<g �<�l�<��<���<��<`   `   خ�<�5�<�5�<��<���<�<���<���<�W�<��<���<��<�E�<3��<��<E�<6��<���<���<X�<��<t��<�<���<`   `   ���<���<���<�w�<e��<�<���<r��<��<�@�<�+�<��<ߨ�<���<��<��<�+�<�@�<��<r��<���<�<F��<�w�<`   `   �K�<	L�<��<�w�<���<��<���<���<���<̕�<1$�<cD�<���<{��<CD�<+$�<���<���<q��<���<��<���<�w�<��<`   `   -�<d=�<)��<��<�a�<�-�<{4�<�V�<�i�<SB�<���<���<���<���<ܷ�<SB�<ci�<�V�<�4�<�-�<Va�<��<J��<d=�<`   `   d=�<ӟ�<�`�<�x�<9��<���< l�<�D�<Z��<�p�<h}�<w
�<�
�<g}�<�p�<l��<E�<l�<u��<X��<�x�<�`�<ɟ�<l=�<`   `   )��<�`�<�2�<�G�<9��< �<���<�9�<t��<��<EU�<&��<5U�<��<���<�9�<���< �<@��<�G�<�2�<�`�<+��<��<`   `   ��<�x�<�G�<}Q�<�y�<���<��<�8�<'9�<��<nS�<lS�<&��<99�<�8�<d�<Ͽ�<�y�<XQ�<�G�<�x�<��<Y��<c��<`   `   �a�<9��<9��<�y�<2i�<�n�<�e�<�B�<f��<D`�<���<D`�<C��<�B�<�e�<�n�<�h�<�y�<u��<9��<la�<��<���<��<`   `   �-�<���< �<���<�n�<	&�<w��<�U�<���<���<���<���<�U�<[��<�%�<�n�<Ͽ�<��<u��<�-�<@��<��<	��<&��<`   `   {4�< l�<���<��<�e�<w��<�(�<Yt�<9��<��<'��<Yt�<�(�<w��<�e�<��<|��< l�<�4�<z�<���<���<���<z�<`   `   �V�<�D�<�9�<�8�<�B�<�U�<Yt�<���<��<��<���<<t�<�U�<�B�<�8�<�9�<E�<�V�<qi�<�y�<+��<��<�y�<�i�<`   `   �i�<Z��<t��<'9�<f��<���<9��<��<��<��<T��<���<7��<'9�<���<Z��<mi�<���<n�<�S�<.f�<�S�<R�<���<`   `   SB�<�p�<��<��<D`�<���<��<��<��<��<���<b`�<&��<���<�p�<[B�<�	�< ��<,1�<<s�<Ws�<Q1�<���<m	�<`   `   ���<h}�<EU�<mS�<���<���<&��<���<T��<���<���<mS�<KU�<h}�<ӷ�<|��<7�<���<�p�<���<�p�<���<h�<|��<`   `   ���<w
�<&��<lS�<D`�<���<Yt�<<t�<���<b`�<mS�<��<�
�<���<M�<��<*�<��<E��<j��<��<�)�<
��<5M�<`   `   ���<�
�<5U�<&��<C��<�U�<�(�<�U�<7��<&��<KU�<�
�<���<A�<��<'��<4<�<�#�<�r�<�#�<@<�<'��<��<A�<`   `   ���<f}�<��<99�<�B�<[��<w��<�B�<'9�<���<h}�<���<A�<�o�<(��<s��<���<���<���<���<���<G��<�o�<0�<`   `   ܷ�<�p�<���<�8�<�e�<�%�<�e�<�8�<���<�p�<ӷ�<M�<��<(��<6�<���<�%�<Α�<I&�<���<��<(��<��<M�<`   `   SB�<l��<�9�<d�<�n�<�n�<��<�9�<Z��<[B�<|��<��<'��<s��<���<��<܎�<���<ܦ�<��<���<��<
��<{��<`   `   ci�<E�<���<Ͽ�<�h�<Ͽ�<|��<E�<mi�<�	�<7�<*�<4<�<���<�%�<܎�<��<܎�<&�<���<*<�<*�<B�<�	�<`   `   �V�<l�< �<�y�<�y�<��< l�<�V�<���< ��<���<��<�#�<���<Α�<���<܎�<��<���<�#�<��<���<���<���<`   `   �4�<u��<?��<XQ�<t��<u��<�4�<qi�<n�<,1�<�p�<E��<�r�<���<I&�<ܦ�<&�<���<s�<E��<�p�<,1�<f�<qi�<`   `   �-�<X��<�G�<�G�<9��<�-�<z�<�y�<�S�<<s�<���<j��<�#�<���<���<��<���<�#�<E��<���<Ws�<�S�<�y�<^�<`   `   Va�<�x�<�2�<�x�<la�<@��<���<+��<.f�<Ws�<�p�<��<A<�<���<��<���<+<�<��<�p�<Ws�<f�<+��<���<@��<`   `   ��<�`�<�`�<��<��<��<���<��<�S�<Q1�<���<�)�<'��<G��<(��<��<*�<���<,1�<�S�<+��<f��<	��<�<`   `   J��<ɟ�<+��<Y��<���<	��<���<�y�<S�<���<h�<
��<��<�o�<��<
��<B�<���<f�<�y�<���<	��<���<Y��<`   `   d=�<l=�<��<c��<��<&��<z�<�i�<���<m	�<|��<5M�<A�<1�<M�<{��<�	�<���<qi�<^�<@��<�<Y��<��<`   `   ��<R�<��<�N�<A��<��<�K�<��<:��<��<1��<���<��<���<J��<��<��<��</L�<��<��<�N�<��<R�<`   `   R�<P��<s��<��<H��<���<T��<��<[��<v��<���<;j�<Lj�<���<Z��<e��<4��<B��<���<[��<�<f��<D��<R�<`   `   ��<s��<��<�<���<���<�}�<rK�<��<�#�<z��<6�<f��<�#�<��<rK�<�}�<���<��<�<޶�<s��<��<��<`   `   �N�<��<�<�p�<���<��<�,�<��<���<��<�.�<�.�<��<���<ġ�<�,�<:��< ��<qp�<�<�<�N�<���<���<`   `   A��<H��<���<���<�C�<I��<G��<���<���<@_�<r��<@_�<|��<���<u��<I��<�C�<���<%��<H��<'��<l��<�V�<l��<`   `   ��<���<���<��<I��<���<d~�<,E�<���<��<��<���<=E�<R~�<���<\��<:��<���<���<��<��<�B�<�B�<ʃ�<`   `   �K�<T��<�}�<�,�<G��<d~�<6�<E��<���<���<���<E��<7�<d~�<P��<�,�<�}�<T��<L�<���<���<f��<Ӝ�<���<`   `   ��<��<qK�<��<���<,E�<E��<��<y��<���<��<3��<=E�<���<ġ�<dK�<4��<��<�r�<�H�<�1�<�1�<�H�<�r�<`   `   :��<[��<��<���<���<���<���<y��<r��<y��<��<���<s��<���<,��<[��<��<R�<+�<Y�<�"�<Y�<�<R�<`   `   ��<v��<�#�<��<@_�<��<���<���<y��<���<��<S_�<��<�#�<Z��<��<�{�<��<z�<�>�<�>�<��<���<�{�<`   `   1��<���<z��<�.�<r��<��<���<��<��<��<b��<�.�<w��<���<K��<Ǌ�<.P�<���<�N�<�p�<IN�<���<[P�<Ǌ�<`   `   ���<;j�<6�<�.�<@_�<���<E��<3��<���<S_�<�.�<6�<Lj�<���<�	�<2E�<�M�<~�<�m�<�m�<��<�M�<&E�<
�<`   `   ��<Lj�<f��<��<|��<=E�<7�<=E�<s��<��<w��<Lj�<��<U��<<��<q�<�3�<o��<�0�<o��<�3�<q�<+��<U��<`   `   ���<���<�#�<���<���<R~�<d~�<���<���<�#�<���<���<U��<���<��<V��<���<�\�<�\�<���<n��<2��<���<D��<`   `   J��<Z��<��<ġ�<u��<���<P��<ġ�<,��<Z��<K��<�	�<<��<��<?�<Q��<"��<��<e��<Q��<
�<��<Y��<�	�<`   `   ��<e��<qK�<�,�<I��<\��<�,�<dK�<[��<��<Ǌ�<2E�<q�<V��<Q��<�9�<M�<+�<�9�<n��<n��<`�<&E�<ˊ�<`   `   ��<4��<�}�<:��<�C�<:��<�}�<4��<��<�{�<.P�<�M�<�3�<���<"��<M�<�u�<M�<&��<���<�3�<�M�<6P�<�{�<`   `   ��<B��<���< ��<���<���<T��<��<R�<��<���<~�<o��<�\�<��<+�<M�<��<�\�<^��<��<���<���<\�<`   `   /L�<���<��<qp�<%��<���<L�<�r�<+�<z�<�N�<�m�<�0�<�\�<e��<�9�<&��<�\�<�0�<�m�<fN�<z�<-�<�r�<`   `   ��<[��<�<�<H��<��<���<�H�<Y�<�>�<�p�<�m�<o��<���<Q��<n��<���<^��<�m�<�p�<�>�<c�<�H�<q��<`   `   ��<�<޶�<�<'��<��<���<�1�<�"�<�>�<IN�<��<�3�<n��<
�<n��<�3�<��<fN�<�>�<�"�<�1�<̜�<��<`   `   �N�<e��<s��<�N�<l��<�B�<f��<�1�<Y�<��<���<�M�<q�<2��<��<`�<�M�<���<z�<c�<�1�<U��<�B�<���<`   `   ��<D��<��<���<�V�<�B�<Ӝ�<�H�<�<���<[P�<'E�<+��<���<Y��<'E�<6P�<���<-�<�H�<̜�<�B�<�V�<���<`   `   R�<R�<��<���<l��<ʃ�<���<�r�<R�<�{�<Ȋ�<
�<U��<D��<�	�<ˊ�<�{�<\�<�r�<q��<��<���<���<��<`   `   ��<d�<�%�<k\�<W��<���<��<�@�<�a�< D�<���<���<z�<���<���< D�<�a�<�@�<��<���<<��<k\�<�%�<d�<`   `   d�<���<s��<
f�<.�<1�<�T�<Gj�<V�<���<��<7��<G��<��<���<V�<aj�<�T�<�0�<.�<f�<o��<���<d�<`   `   �%�<s��<�6�<y��<��<��<���<���<YI�<��<a�<)��<�`�<��<nI�<���<��<��<-��<y��<~6�<s��<�%�<���<`   `   k\�<
f�<y��<G��<+x�<�a�<\3�<���<�(�<"�<���<���<1�<�(�<���<V3�<�a�<2x�<.��<u��<f�<g\�<���<��<`   `   W��<.�<��<+x�<�D�<��<���<6��<
��<���<8��<���<���<6��<���<��<�D�<+x�<8��<.�<G��<!9�<1��<!9�<`   `   ���<1�<��<�a�<��<��<���<��<s�<P��<I��<s�<��<���<��<��<�a�<��<�0�<���<���<#�<�<���<`   `   ��<�T�<���<\3�<���<���<ٹ�<�l�<J��<P�<O��<�l�<ѹ�<���<���<\3�<��<�T�<��</�<{a�<�(�<�a�</�<`   `   �@�<Gj�<���<���<6��<��<�l�<}��<�<�<v��<�l�<��<=��<���<���<aj�<�@�</A�<���<$�<$�<���<GA�<`   `   �a�<V�<YI�<�(�<
��<s�<J��<�<T�<�<W��<s�<���<�(�<sI�<V�<�a�<��<���<�N�<$�<�N�<���<��<`   `    D�<���<��<"�<���<O��<P�<�<�<J�<I��<���<1�<���<���<�C�<H��<d��<y�<�4�<�4�<4y�<X��<.��<`   `   ���<��<a�<���<8��<I��<O��<v��<W��<I��<7��<���<�`�<��<���<8Q�<���<�s�<�)�<��<�)�<�s�<���<8Q�<`   `   ���<7��<)��<���<���<s�<�l�<�l�<s�<���<���<%��<F��<|��<:��<�Y�<��<���<Ѱ�<��<���<��<�Y�<P��<`   `   z�<F��<�`�<1�<���<��<ѹ�<��<���<1�<�`�<F��<n�<@7�<	K�<>�<��<P��<O��<P��<��<>�<�J�<@7�<`   `   ���<��<��<�(�<6��<���<���<=��<�(�<���<��<|��<@7�< ��<���<k��<���<��<���<���<��<���<���<17�<`   `   ���<���<nI�<���<���<��<���<���<sI�<���<���<:��<	K�<���<+�<T�<�`�<�b�<�`�<T�<�*�<���<%K�<:��<`   `    D�<V�<���<V3�<��<��<\3�<���<V�<�C�<8Q�<�Y�<>�<k��<T�<��<���<r��<���<+T�<��<>�<�Y�<?Q�<`   `   �a�<aj�<��<�a�<�D�<�a�<��<aj�<�a�<H��<���<��<��<���<�`�<���<��<���<�`�<���<��<��<���<H��<`   `   �@�<�T�<��<2x�<+x�<��<�T�<�@�<��<d��<�s�<���<P��<��<�b�<r��<���<�b�<���<A��<���<�s�<X��<��<`   `   ��<�0�<-��<.��<7��<�0�<��</A�<���<y�<�)�<Ѱ�<O��<���<�`�<���<�`�<���<w��<Ѱ�<�)�<y�<���</A�<`   `   ���<.�<y��<u��<.�<���</�<���<�N�<�4�<��<��<P��<���<T�<+T�<���<A��<Ѱ�<��<�4�<�N�<���<(�<`   `   <��<f�<~6�<f�<G��<���<{a�<$�<$�<�4�<�)�<���<��<��<�*�<��<��<���<�)�<�4�<�#�<$�<�a�<���<`   `   k\�<o��<s��<g\�<!9�<#�<�(�<$�<�N�<4y�<�s�<��<>�<���<���<>�<��<�s�<y�<�N�<$�<�(�<�<(9�<`   `   �%�<���<�%�<���<1��<�<�a�<���<���<X��<���<�Y�<�J�<���<%K�<�Y�<���<X��<���<���<�a�<�<6��<���<`   `   d�<d�<���<��<!9�<���</�<HA�<��<.��<8Q�<P��<A7�<17�<:��<?Q�<H��<��</A�<(�<���<(9�<���<���<`   `   ���<@'�<ƣ�<gb�<zY�<�q�<�<���<��<�f�<��<�B�<�]�<�B�<��<�f�<��<���<ʖ�<�q�<rY�<gb�<ʣ�<@'�<`   `   @'�<W��<$��<z��<A�<���<�O�<%��<\��<N��<Ԁ�<&��<2��<݀�<A��<U��<3��<�O�<���< A�<���<+��<M��<8'�<`   `   ƣ�<$��<r��<Ӳ�<��<�z�<�@�<���<��<r	�<���<���<r��<r	�<�<���<�@�<�z�<)��<Ҳ�<_��<$��<٣�<�K�<`   `   gb�<z��<Ҳ�<F��<��<�=�<�&�<Ż�<���<���<#1�<,1�<���<���<���<�&�<>�<��<8��<ٲ�<���<_b�<���<��<`   `   yY�<A�<��<��<u��<���<���<�H�<^Y�<���<5�<���<ZY�<�H�<���<���<l��<��<��<A�<uY�<��<��<��<`   `   �q�<���<�z�<�=�<���<�#�<$��<Y�<9�<���<���<9�<�Y�<*��<�#�<���<>�<�z�<���<�q�<���<%��<��<���<`   `   �<�O�<�@�<�&�<���<$��<)��<M��<q��<���<���<M��<��<$��<���<�&�<�@�<�O�<ؖ�<�h�<���<�y�<��<�h�<`   `   ���<%��<���<Ż�<�H�<Y�<M��<���<{J�<tJ�<���<S��<�Y�<�H�<���<���<3��<~��<`�<��<�	�<�	�<��<n�<`   `   ��<\��<��<���<^Y�<9�<q��<{J�<���<{J�<t��<9�<XY�<���<��<[��<��<���<>�<[e�<���<[e�<;�<���<`   `   �f�<N��<r	�<���<���<���<���<tJ�<{J�<���<���<���<���<y	�<A��<�f�<���<���<���<E�< E�<���<���<���<`   `   ��<Ԁ�<���<#1�<5�<���<���<���<t��<���<!5�<#1�<t��<Ӏ�<*��<�+�<���<���<�z�<���<�z�<���<���<�+�<`   `   �B�<&��<���<,1�<���<9�<M��<S��<9�<���<#1�<���<1��<�B�<�D�<�0�<�z�<c��<x�<��<p��<�z�<�0�<�D�<`   `   �]�<1��<r��<���<ZY�<�Y�<��<�Y�<XY�<���<t��<1��<�]�<�M�<L��<_��<}�<~��<ӳ�<~��<�<_��<I��<�M�<`   `   �B�<܀�<r	�<���<�H�<)��<$��<�H�<���<y	�<Ӏ�<�B�<�M�<8��<i(�<v��<8��<#��<��<*��<���<v(�<.��<�M�<`   `   ��<A��<�<���<���<�#�<���<���<��<A��<*��<�D�<L��<i(�<�z�<K}�<���<mֿ<���<K}�<hz�<i(�<b��<�D�<`   `   �f�<U��<���<�&�<���<���<�&�<���<[��<�f�<�+�<�0�<_��<v��<K}�<}�<�8�<�8�<o�<X}�<���<T��<�0�<�+�<`   `   ��<3��<�@�<>�<l��<>�<�@�<3��<��<���<���<�z�<~�<8��<���<�8�<sQ�<�8�<���<8��<|�<�z�<���<���<`   `   ���<�O�<�z�<��<��<�z�<�O�<~��<���<���<���<c��<~��<#��<mֿ<�8�<�8�<zֿ<��<s��<p��<���<���<���<`   `   ʖ�<���<)��<8��<��<���<ؖ�<`�<?�<���<�z�<y�<ӳ�<��<���<o�<���<��<��<y�<�z�<���<P�<`�<`   `   �q�< A�<Ҳ�<ٲ�<A�<�q�<�h�<��<[e�<E�<���<��<~��<*��<K}�<X}�<8��<s��<y�<��< E�<Te�<��<�h�<`   `   rY�<���<^��<���<uY�<���<���<�	�<���< E�<�z�<p��<�<���<hz�<���<|�<p��<�z�< E�<���<�	�<���<���<`   `   gb�<+��<$��<_b�<��<%��<�y�<�	�<[e�<���<���<�z�<_��<v(�<i(�<T��<�z�<���<���<Te�<�	�<�y�<��<��<`   `   ʣ�<M��<٣�<���<��<��<��<��<;�<���<���<�0�<I��<.��<b��<�0�<���<���<P�<��<���<��<���<���<`   `   @'�<8'�<�K�<��<��<���<�h�<n�<���<���<�+�<�D�<�M�<�M�<�D�<�+�<���<���<`�<�h�<���<��<���<�K�<`   `   �<2��<��<�/�<�w�<�i�<���<���<W��<�}�<��<�3�<���<�3�<��<�}�<f��<���<���<�i�<�w�<�/�<ۨ�<2��<`   `   2��<�,�<��<Y��<^�<��<�E�<���<���<���<���<���<���<���<���<���<��<�E�<��<^�<\��<'��<�,�<&��<`   `   ��<��<���<�Y�<��<v�<���<�]�<It�<�U�<�1�<p �<�1�<�U�<Yt�<�]�<���<u�<.��<�Y�<���<��<���<]Z�<`   `   �/�<Y��<�Y�<���<�m�<؞�<�W�<t��<E�<���<��<��<���<qE�<s��<�W�<מ�<�m�<���<�Y�<\��<�/�<�,�<�,�<`   `   �w�<^�<��<�m�<|��<���<�&�<���<���<�w�<���<�w�<���<���<}&�<���<���<�m�<��<^�<�w�<��<��<��<`   `   �i�<��<u�<؞�<���<yX�<{�<��<�H�<���<���<�H�<��<��<xX�<���<מ�<��<��<�i�<N�<؜�<М�<N�<`   `   ���<�E�<���<�W�<�&�<{�<�"�<�3�<I`�<o��<a`�<�3�<�"�<{�<�&�<�W�<���<�E�<���<�~�<y��<j��<���<�~�<`   `   ���<���<�]�<t��<���<��<�3�<F<�<0A�<!A�<<<�<4�<��<q��<s��<�]�<��<���<��<͡�<�>�<�>�<ơ�<��<`   `   W��<���<It�<E�<���<�H�<I`�<0A�<9��<0A�<A`�<�H�<���<E�<:t�<���<d��<H4�<��<;׮<�g�<;׮<"��<H4�<`   `   �}�<���<�U�<���<�w�<���<n��<!A�<0A�<���<���<�w�<���<�U�<���<�}�<7�<��<C��<�\�<�\�<C��<��<7�<`   `   ��<���<�1�<��<���<���<a`�<<<�<A`�<���<���<��<�1�<���<��<���<.�<8��<�ʘ<QƖ<�ʘ<8��<.�<���<`   `   �3�<���<o �<��<�w�<�H�<�3�<4�<�H�<�w�<��< �<���<~3�<8ͮ<X�<+�<c��<��<��<f��<	+�<�W�<9ͮ<`   `   ���<���<�1�<���<���<��<�"�<��<���<���<�1�<���<��<H�<_�<⎑<:=�<]`}<�x<]`}<6=�<⎑<f�<H�<`   `   �3�<���<�U�<qE�<���<��<{�<q��<E�<�U�<���<~3�<H�<���<L��<}��<T�k<�}`<�}`<U�k<���<M��<x��<zH�<`   `   ��<���<Xt�<s��<}&�<xX�<�&�<s��<:t�<���<��<8ͮ<_�<L��<9<}<��b<)�P<�vJ<'�P<��b<1<}<L��<l�<8ͮ<`   `   �}�<���<�]�<�W�<���<���<�W�<�]�<���<�}�<���<X�<⎑<}��<��b<�/K<��><��><�/K<��b<���<ݎ�<�W�<���<`   `   f��<��<���<מ�<���<מ�<���<��<d��<7�<.�<+�<:=�<T�k<)�P<��><48<��><'�P<T�k<<=�<+�<.�<7�<`   `   ���<�E�<u�<�m�<�m�<��<�E�<���<H4�<��<8��<c��<]`}<�}`<�vJ<��><��><�vJ<�}`<S`}<f��<B��<��<:4�<`   `   ���<��<-��<���<��<��<���<��<��<D��<�ʘ<��<�x<�}`<(�P<�/K<'�P<�}`<�x<��<zʘ<D��<0��<��<`   `   �i�<^�<�Y�<�Y�<^�<�i�<�~�<͡�<<׮<�\�<QƖ<��<]`}<V�k<��b<��b<T�k<T`}<��<[Ɩ<�\�<-׮<ơ�<�~�<`   `   �w�<\��<���<\��<�w�<N�<y��<�>�<�g�<�\�<�ʘ<f��<7=�<���<2<}<���<<=�<f��<zʘ<�\�<�g�<�>�<o��<N�<`   `   �/�<'��<��<�/�<��<؜�<k��<�>�<<׮<D��<8��<	+�<⎑<N��<L��<ݎ�<+�<B��<D��<-׮<�>�<|��<М�<���<`   `   ۨ�<�,�<���<�,�<��<ќ�<���<ơ�<"��<��<.�<�W�<f�<y��<l�<�W�<.�<��<0��<ơ�<o��<М�<2��<�,�<`   `   2��<&��<]Z�<�,�<��<N�<�~�<��<H4�<7�<���<9ͮ<H�<zH�<8ͮ<���<7�<:4�<��<�~�<N�<���<�,�<nZ�<`   `   ZX�<Y��<���<���<^ʹ<�8�<2�<�<G�<��<j\�<G��<!�<G��<S\�<��<n�<�<�1�<�8�<�ʹ<���<o��<Y��<`   `   Y��<�V�<w��<T3�<�(�<�(�<�<�+�<�٧<�ע<��<h̜<e̜<�<�ע<y٧<�+�<"�<�(�<�(�<K3�<���<V�<J��<`   `   ���<w��<�N�<��<�E�<B˽<r�<{X�<�ط<ku�<�<��<췳<ku�<�ط<{X�<r�<B˽<�E�<��<�N�<w��<���<�Ļ<`   `   ���<T3�<��<c��<�u�<�I�<�=�<�^�<���<J�<���<��<J�<���<�^�<�=�<tI�<nu�<s��<��<K3�<���<�ͷ<�ͷ<`   `   ^ʹ<�(�<�E�<�u�<�(�<���<_��<���<�{�<���<w��<���<�{�<���<6��<���<)�<�u�<�E�<�(�<vʹ<`ر<�ϰ<`ر<`   `   �8�<�(�<B˽<�I�<���<���<���<U��<�S�<+�<+�<�S�<R��<ï�<���<���<tI�<[˽<�(�<�8�<��<���<���<��<`   `   2�<�<r�<�=�<_��<���<k��<�y�<~��<qH�<���<�y�<R��<���<p��<�=�<r�<�<2�<5�<�V�<�g�<�V�<5�<`   `   �<�+�<{X�<�^�<���<U��<�y�<=b�<vS�<aS�<4b�<�y�<R��<e��<�^�<�X�<�+�<	�<�<�$�<�Q�<�Q�<�$�<�<`   `   G�<�٧<�ط<���<�{�<�S�<~��<vS�<��<vS�<k��<�S�<�{�<���<�ط<�٧<h�<�0�<5t<7�b<Dy\<7�b<\t<�0�<`   `   ��<�ע<ku�<J�<���<
+�<qH�<aS�<vS�<�H�<+�<~��<J�<�u�<�ע<��<�t<'@P<"�4<.&<&<�4<"@P<�t<`   `   i\�<��<�<���<w��<+�<���<4b�<k��<+�<���<���<ܷ�<��<k\�<GG]<OF.<U*<H�;���;�H�;U*<0F.<GG]<`   `   G��<h̜<��<��<���<�S�<�y�<�y�<�S�<~��<���<�<d̜<8��<h�K<G<�g�;dB[;��;R�;B[;?h�;B<N�K<`   `    �<d̜<췳<J�<�{�<Q��<Q��<Q��<�{�<J�<ܷ�<d̜<3�<a=B<�~�;W�|;��:�~Ӻ9��~Ӻ��:X�|;�~�;b=B<`   `   G��<�<ju�<���<���<ï�<���<e��<���<�u�<��<8��<a=B<?J�;�<9;v����;��\�ǻ�ǻp;�����'<9;4J�;h=B<`   `   S\�<�ע<�ط<�^�<6��<���<p��<�^�<�ط<�ע<k\�<h�K<�~�;�<9;����}���y���3����|���0����<9;�~�;h�K<`   `   ��<y٧<{X�<�=�<���<���<�=�<�X�<�٧<��<GG]<H<X�|;u���}���X�k�:�F�:�7��������s�|;B<YG]<`   `   m�<�+�<r�<sI�<)�<sI�<r�<�+�<h�<�t<OF.<�g�;��:�;��x��j�:�hK�j�:����;��c�:�g�;CF.<�t<`   `   �<"�<B˽<mu�<�u�<[˽<�<	�<�0�<(@P<U*<eB[;�~Ӻ[�ǻ�3�F�:�j�:��3��ǻM~ӺB[;g*<"@P<�0�<`   `   �1�<�(�<�E�<s��<�E�<�(�<2�<�<6t<#�4<H�;��;9��ǻ���7����ǻ�9���;H�;#�4<dt<�<`   `   �8�<�(�<��<��<�(�<�8�<5�<�$�<7�b</&<���;T�;�~Ӻo;��|��������;��L~Ӻ��;���;&<�b<�$�<Q�<`   `   �ʹ<K3�<�N�<K3�<vʹ<��<�V�<�Q�<Ey\<&<�H�; B[;��:����,�������h�: B[;H�;&<�y\<�Q�<rV�<��<`   `   ���<���<w��<���<`ر<���<�g�<�Q�<7�b<�4<U*<@h�;[�|;)<9;�<9;u�|;�g�;h*<#�4<�b<�Q�<�g�<���<Bر<`   `   o��<V�<���<�ͷ<�ϰ<���<�V�<�$�<\t<#@P<1F.<C<�~�;6J�;�~�;C<CF.<#@P<et<�$�<rV�<���<�ϰ<�ͷ<`   `   Y��<J��<�Ļ<�ͷ<`ر<��<5�<�<�0�<�t<GG]<N�K<b=B<i=B<i�K<ZG]<�t<�0�<�<R�<��<Bر<�ͷ<�Ļ<`   `   Uc�<(��<��<�k�<�ח<��<<�q<�J<� <.��;�;k�};��];k�};��;.��;& <�J<��q<��<�ח<�k�<���<(��<`   `   (��<蘬<i��<,�<�d�<\m�<R1�<��z<r�_<N�F<��3<�8)<�8)<Ƽ3<��F<>�_<Z�z<x1�<~m�<�d�<�<���<올<��<`   `   ��<i��<�Y�<ZQ�<]�<��<�M�<6Y�<�<W}�<��<FH�<��<W}�<��<6Y�<�M�<��<c�<ZQ�<�Y�<i��<'��<���<`   `   �k�<,�<ZQ�<�g�<���<�8�<�U�<3�<�y�<4�<B��<I��<'�<�y�<"3�<�U�<j8�<[��<	h�<zQ�<�<�k�<���<���<`   `   �ח<�d�<]�<���<d�<��<��<��<��<!�<+�<!�<��<��<r�<��<��<���<�<�d�<�ח<�v�<��<�v�<`   `   ��<\m�<��<�8�<��<�{�<���<K��<��<��<x��<��<=��<���<�{�<��<j8�<��<~m�<��<�!�<ưx<Ͱx<�!�<`   `   ;�q<R1�<�M�<�U�<��<���<�y�<�u�<K��<��<l��<�u�<qy�<���<��<�U�<�M�<R1�<�q<WQT<I�@<L�9<�@<WQT<`   `   �J<��z<6Y�<3�<��<K��<�u�<F�<=��<#��<F�<�u�<=��<ے�<"3�<VY�<Y�z<xJ<�i<Q�;A2�;�2�;Q�;�i<`   `   � <q�_<�<�y�<��<��<K��<=��<C��<=��<,��<��<��<�y�<��<q�_< <���;�B;y�o:�_F9z�o:�B;���;`   `   -��;M�F<W}�<4�<!�<��<��<#��<=��<��<x��<� �<'�<w}�<��F<��;er ;��
ʫ����ݣ滔ʫ�����s ;`   `   �;��3<��<B��<+�<x��<k��<F�<,��<x��<Z�<B��<��<��3<��;��Q���׻�x;�ڕp�=���i�p��x;�\�׻��Q�`   `   h�};�8)<EH�<I��<!�<��<�u�<�u�<��<� �<B��<fH�<�8)<�};��U��+�&�������ʼ=�ʼ�������+���U�`   `   ��];�8)<��<'�<��<=��<qy�<=��<��<'�<��<�8)<��];y���QzV�ځ���R��������S�ځ��zV�x���`   `   h�};Ƽ3<W}�<�y�<��<���<���<ے�<�y�<w}�<��3<�};y���Fxe�����` �G}/�6}/�` ���,��?xe�D���`   `   ��;��F<��<"3�<r�<�{�<��<"3�<��<��F<��;��U�PzV���%�
��X.�
kF�I�N�.kF��X.��
���qzV���U�`   `   -��;>�_<5Y�<�U�<��<��<�U�<VY�<q�_<��;��Q��+�ځ�����X.���N��$`�|$`��N�Y.���́���+���Q�`   `   % <Y�z<�M�<i8�<��<i8�<�M�<Y�z< <fr ;��׻&����R�` �
kF��$`�FAi��$`�kF�` ��R�&�����׻gr ;`   `   �J<x1�<��<[��<���<��<R1�<xJ<���;���x;������G}/�I�N�|$`��$`�W�N�5}/�������x;����4��;`   `   ��q<~m�<c�<	h�<�<~m�<�q<�i<�B;	ʫ�ٕp��ʼ���5}/�.kF��N�kF�5}/�Ё��ʼ��p�	ʫ���B;�i<`   `   ��<�d�<ZQ�<zQ�<�d�<��<WQT<Q�;��o:���<���=�ʼ��` ��X.�Y.�` ����ʼ5���ۣ�L�o:Q�;�QT<`   `   �ח<�<�Y�<�<�ח<�!�<J�@<B2�;!`F9ۣ�h�p����S����
����R������p�ۣ�
xF9B2�;��@<�!�<`   `   �k�<���<i��<�k�<�v�<ưx<L�9<�2�;��o:�ʫ��x;� ���ځ��,����́��%����x;�	ʫ�O�o:C2�;��9<Ͱx<�v�<`   `   ���<올<'��<���<��<Ͱx<�@<Q�;�B;���Z�׻�+�zV�>xe�qzV��+���׻�����B;Q�;��@<Ͱx<�<���<`   `   (��<��<���<���<�v�<�!�<WQT<�i<���;�s ;��Q��U�w���B�����U���Q�ir ;5��;�i<�QT<�!�<�v�<���<���<`   `   ���<R�<Տ<Pz�<��X<�l!<xY�;vk:u��_,���X�F7��59��F7����X�_,��s��vk:�W�;�l!<s�X<Pz�<�ԏ<R�<`   `   R�<��<�ߎ<D��<Ɉl<{lF<w�<'��;��0;�y���C1��䂻P傻kC1�n����0;E��;ӹ<�lF<f�l< ��<�ߎ<��<@�<`   `   Տ<�ߎ<���<F}�<֒�<��n<4JT<��5<Z�<��;"��;?��;r��;��;9�<��5<HJT<��n<Ӓ�<E}�<���<�ߎ<$Տ<R�<`   `   Pz�<D��<E}�<�y�<%�<�ˊ<�{�<�N�<N=s<� h<:�a<A�a<| h<=s<�N�<�{�<ˊ<�~�<�y�<m}�< ��<?z�<�*<�*<`   `   ��X<Ɉl<֒�<%�<;p�<$��<ѽ�<ɚ�<�,�<+y�<!)�<+y�<�,�<ɚ�<u��<$��<�p�<%�<z��<Ɉl<1�X<��K<G<��K<`   `   �l!<zlF<��n<�ˊ<$��<n��<_�<R��<��<�!�<�!�<�<:��<��<���<�<ˊ<��n<�lF<�l!<U<��;7��;�<`   `   wY�;v�<3JT<�{�<ѽ�<_�<��<{��<���<���<���<{��<��<_�<ս�<�{�<UJT<v�<�X�;��/;!�/:�]�^�/:��/;`   `   vk:&��;��5<�N�<ɚ�<Q��<{��<��<)�<�<
��<���<:��<���<�N�<D�5<D��;�sk:s�u�T�z;�3;�*��u�`   `   u����0;Z�<N=s<�,�<��<���<)�<R��<)�<o��<��<�,�<N=s<��<��0;�s���x1��z��*������*��bz���x1�`   `   _,��y����;� h<+y�<�!�<���<�<)�<ӯ�<�!�<�x�<{ h<<�;;n���,�7����ռ�M�p����M���ռ����`   `   ��X��C1� ��;9�a< )�<�!�<���<
��<o��<�!�<V)�<9�a<���;�C1���X���ȼ�0��7�СP�ɦY���P��7��0���ȼ`   `   F7���䂻=��;@�a<+y�<�<{��<���<��<�x�<9�a<���;R傻X7����|y1���e�߆��ᑽ�ᑽ߆�w�e�wy1���`   `   59��Q傻q��;{ h<�,�<9��<��<9��<�,�<{ h<���;R傻9��)��a+G�u���c�2)��q���2)��h�u���O+G�)��`   `   F7��nC1���;=s<ɚ�<��<_�<���<M=s<<�;�C1�X7��)����N��m��^���_�ν\e޽Oe޽Q�νf����m����N���`   `   ��X�2n��8�<�N�<u��<���<ս�<�N�<��<:n����X���a+G��m��%丽׈ݽ���H|�����׈ݽ丽�m��q+G���`   `   _,���0;��5<�{�<#��<�<�{�<D�5<��0;�,���ȼ|y1�u���^���׈ݽ.-��q��i�� -���ݽf���o���wy1���ȼ`   `   �s��D��;GJT<ˊ<�p�<ˊ<UJT<D��;�s��7����0���e�c�_�ν���q��{��q�����_�ν`򠽓�e��0�6���`   `   vk:ҹ<��n<�~�<%�<��n<v�<�sk:�x1��ռ�7�߆�2)��\e޽H|��i��q��S|��Oe޽,)��߆��7���ռ�x1�`   `   �W�;�lF<Ӓ�<�y�<y��<�lF<�X�;r�u��z���M�СP��ᑽq���Oe޽��� -�����Oe޽�����ᑽ��P��M�yz��q�u�`   `   �l!<e�l<E}�<l}�<Ɉl<�l!<��/;S�*��o�ɦY��ᑽ2)��Q�ν׈ݽ�ݽ_�ν,)���ᑽǦY���;*��*�m�/;`   `   r�X< ��<���< ��<1�X<U<'�/:z;���������P�߆�h�f���丽f���`�߆���P���R���z;��/:U<`   `   Pz�<�ߎ<�ߎ<?z�<��K<��;]�2;�*���M��7�w�e�u����m���m��o�����e��7��M�;*��z;�� �7��;��K<`   `   �ԏ<��<$Տ<�*<G<7��;g�/:)�az����ռ�0�wy1�O+G���N�q+G�wy1��0���ռyz��)��/:7��;nG<�*<`   `   R�<@�<R�<�*<��K<�<��/;�u��x1�������ȼ��)�������ȼ6����x1�p�u�n�/;U<��K<�*<y�<`   `   J�}<зt<+7X<�K&<���;������2ㅼ�UѼ�R�!l,��jA��H��jA�@l,��R�<UѼ2ㅼm��������;�K&<�6X<зt<`   `   зt<G+j<��S<}�.<:��;K�Q;���{ ���c��Y���{¼��ռ��ռ�{¼�Y����c��{ ����|�Q;S��;�.<ܘS<i+j<��t<`   `   +7X<��S</�I<�S7<\�<Ah�;���;�U�9��G��Oǻ�c��T��c��Oǻ��G��U�9��;Ah�;C�<�S7<9�I<��S<*7X<��Y<`   `   �K&<}�.<�S7<'O<<#:<��.<�<�9<���;���;���;���;��;@��;d:<��<8�.<�":<�O<<"T7<�.<^K&<. !< !<`   `   �;9��;\�<#:<�}R<�wa<�+g<��e<��a<�>]< �[<�>]<�a<��e<�*g<�wa<�~R<#:<w�<9��;���;{��;�w�;{��;`   `   ��I�Q;@h�;��.<�wa<�<ր�<2��<�v�<�m�<�m�<�v�<��<��<R�<Wwa<7�.<�h�;y�Q;*� �F�����Y�����F�`   `   ����������;�<�+g<ր�<H7�<L}�<�i�<K�<�i�<L}�<67�<ր�<�+g<�</��;���V���c�N�A ������ ��c�N�`   `   3ㅼ{ �sU�9�9<��e<2��<L}�<2��<~�<_�<2��<�}�<��<4�e<c:<�`�9�{ �Dㅼ#eżL ��yW�aW�; ��ież`   `   �UѼ��c���G����;��a<�v�<�i�<~�<.��<~�<ai�<�v�<C�a<���;��G���c�KUѼv#��>�4Y�@�b�4Y���>�v#�`   `   �R��Y���Oǻ���;�>]<�m�<K�<_�<~�<��<�m�<�>]<��;!Oǻ�Y���R���L�����l���ئ�٦��l�� �����L�`   `   !l,��{¼�c����;��[<�m�<�i�<2��<`i�<�m�<q�[<���;�c��{¼7l,�	I~������+ʽ^���@���+ʽ����	I~�`   `   �jA���ռ�T����;�>]<�v�<L}�<�}�<�v�<�>]<���;9T���ռ�jA�4��ƽ�����D��������D�����ƽ"4��`   `   �H���ռ�c���;�a<��<57�<��<B�a<��;�c���ռe�H�������ڽ{����'���:�6/A���:���'�{����ڽ����`   `   �jA��{¼�Oǻ>��;��e<
��<ր�<4�e<���;!Oǻ�{¼�jA������:�T2��X9�_>U���d���d�U>U��X9�[2��:�z���`   `   @l,��Y����G�c:<�*g<R�<�+g<c:<��G��Y��7l,�4����ڽT2��?��d��t}�G��u}��d�q�?�T2���ڽ4��`   `   �R���c�jU�9��<�wa<Wwa<�<~`�9��c��R�	I~�ƽ{���X9��d��(�����������(���d��X9�w��ƽ	I~�`   `   <UѼ�{ ���;7�.<�~R<7�.</��;�{ �KUѼ��L�����������'�_>U��t}������������t}�_>U�~�'�����������L�`   `   2ㅼ��?h�;�":<#:<�h�;���Dㅼu#�����+ʽ�D���:���d�G����������G����d���:��D��+ʽ ����#�`   `   n���y�Q;B�<�O<<v�<y�Q;V���#eż�>��l��^�὿��6/A���d�u}��(���t}���d�C/A����Q�Ὧl���>�#eż`   `   ��S��;�S7<"T7<8��;(�c�N�L ��4Y��ئ�������:�U>U��d��d�_>U���:�����٦�4Y�; ����N�`   `   ���;�.<8�I<�.<���;�F�A ��yW�?�b�٦�@�ὰD���'��X9�q�?��X9�~�'��D�Q��٦��b�yW�� ���F�`   `   �K&<ܘS<��S<^K&<{��;�������`W�4Y��l���+ʽ����{��[2�T2�w�������+ʽ�l��4Y�yW�΅��X������;`   `   �6X<i+j<*7X<. !<�w�;X���� ��: ����>� �������ƽ��ڽ�:���ڽƽ���� ����>�: ��� ��X����x�;. !<`   `   зt<��t<��Y< !<{��;��F�b�N�ieżu#���L�	I~�"4������z���4��	I~���L��#�"eż��N��F����;. !<�Y<`   `   �A6<)�'<�c�;��);B�����k�3lڼ@)(��h�����l�����z7ǽ����l������h�A)(��lڼ��k�R�����);�b�;)�'<`   `   )�'</z<t�;��V;=���b����W��(��ȇA���_���o�	�o���_���A�8�����~��b�:����V;�t�;]z<�'<`   `   �c�;t�;2S�;u~;��a:�Z������m�
ݧ�+Ҽ�������a��+Ҽ5ݧ���m�}���Z���a:u~;bS�;t�;�c�;/�;`   `   ��);��V;u~;��;O;e;�z;I�n�O@F��Y�����/��8��-��yZ���=F�kxn�#x;R9e;a�;�v~;��V;:�);�a;�`;`   `   B���>����a:O;e;��;s�;���;���;���;QO�;-�;QO�;۹�;���;���;s�;'!�;N;e;�sa:?������һ���һ`   `   ��k��b��Z��z;s�;Io"<��G<�]<��h<km<km<��h<��]<&�G<�o"<r�;!x;Z�b���k�߾��eH��MH������`   `   4lڼ������g�n����;��G<wx�<H�<��<̍�<��<H�<ix�<��G<���;��n�k�����ylڼmj��o!�p�(��o!�mj�`   `   A)(�W�Ἦ�m�Q@F����;�]<H�<h�<�u�<�u�< h�<��<��]<���;�=F�N�m����I)(��[��7��z���k����7���[�`   `   �h�(��
ݧ��Y�����;��h<��<�u�<'��<�u�<W�<��h<S��;�Y���ݧ�(���h��/��s꺽�/ѽ�ٽ�/ѽd꺽�/��`   `   ���ɇA�+Ҽ���PO�;km<̍�<�u�<�u�<��<km<QN�;.���Ҽ��A����b�ȽϏ��s���ʘ�~��ɏ��L�Ƚ`   `   �l����_����0��-�;km<��<h�<W�<km<�-�;0�����_��l��%����&�;���P��_X���P�&�;���%��`   `   �����o�����8��OO�;��h<H�<��<��h<QN�;0������
�o����� �%�8�M�d�Ѳ��,o��2o��Բ��B�d�"�8��`   `   z7ǽ	�o�a��.��ٹ�;��]<ix�<��]<R��;.�����
�o�k7ǽrZ���K��}��.�)���T+��)���/򛾌}����K�rZ�`   `   �����_�+Ҽ{Z�����;%�G<��G<���;�Y���Ҽ��_����rZ�6�R����1ᬾ��Ǿ�8׾�8׾{�Ǿ4ᬾ���3�R�mZ�`   `   �l����A�5ݧ��=F����;�o"<���;�=F��ݧ���A��l��� ���K����|���r�־l�u9��w�r�־s��������K�� �`   `   ���8����m��xn�s�;r�;��n�N�m�(�����%��%�8��}��1ᬾr�־$
��&I�$I�
��v�־4ᬾ�}��"�8�&��`   `   �h����~�� x;&!�;x;l����Ἵh�b�Ƚ��M�d�.򛾁�Ǿl�&I�{�&I�l��Ǿ,�M�d���b�Ƚ`   `   A)(�~���Z�P9e;K;e;	Z����I)(��/��Ϗ��%�;�в��)����8׾u9��$I�&I�z9���8׾&���Բ��&�;�ɏ���/��`   `   �lڼb��a:`�;�sa:b�ylڼ�[�s꺽s����P�,o��T+���8׾w�
��l�8׾\+��,o����P�s��p꺽�[�`   `   ��k�<��u~;�v~;@����k�mj��7���/ѽ��_X�2o��)���{�Ǿr�־v�־��Ǿ&���,o���_X�ʘ��/ѽ�7��Pj�`   `   R�����V;aS�;��V;���߾���o!�z����ٽʘ���P�Բ��/�4ᬾs���4ᬾ,�Բ����P�ʘ��ٽz����o!�߾��`   `   ��);�t�;t�;9�);�һdH��o�(�k����/ѽ~��%�;�A�d��}���������}��M�d�&�;�s���/ѽz���S�(�MH���һ`   `   �b�;]z<�c�;�a;��MH���o!��7��c꺽ɏ����"�8���K�3�R���K�"�8���ɏ��p꺽�7���o!�MH��K軳a;`   `   )�'<�'</�;�`;�һ����mj��[��/��K�Ƚ%���rZ�mZ�� �&��b�Ƚ�/���[�Pj�߾���һ�a;��;`   `   �u�;+̑;K�9�
㻧��xO�ƠT�����E`̽����H>%�Ϊ*�H>%�$����"`̽�����T�xO����
�K7�9+̑;`   `   +̑;��<;�����Ż@�g���̼�����]��N��x���ǽv&ս�&ս�ǽx���N����]�e����̼ȶg���Ż��h�<;�ˑ;`   `   K�9������sY��#$&�zd����ͼ�l�p^4��V��m�=u��m��V��^4��l���ͼzd��^$&�tY��3�����8H�9ò:`   `   �
㻕�ŻsY�����Ɯ׻�����S��m���Ӵ�^Ӽ�����㼒ӼԴ�gm��m�S�{��՝׻~����X����Ż>�8�������`   `   ���A�g�#$&�Ɯ׻�΄�+�:�tR>��z�h���@Ȼk1ջ�@Ȼ�f���z�W>�,�:�	̄�ǜ׻M%&�A�g�Q��`^��#��`^��`   `   xO���̼zd�����,�:��J�:gך;W��;��;��;	��;���;���;\ؚ;
P�:K�:�{��Gd����̼�O�7���,���,��6�`   `   ƠT������ͼ��S�uR>�gך;��$<-\<̽y<Kx�<��y<-\<��$<fך;S>���S���ͼ����T��ǁ�@���:[��X����ǁ�`   `   ������]��l��m���z�V��;-\<�j�<
�<�	�<�j�<�\<���;?�z�gm���l���]�����5��^�޽��ｕ��W�޽+5��`   `   E`̽�N��p^4��Ӵ�h����;̽y<
�<���<
�<A�y<��;7f���Ӵ��^4��N��'`̽9I��s��h0�'�6��h0��s�9I�`   `   ���x���V�^Ӽ�@Ȼ��;Kx�<�	�<
�<�x�<��;�AȻ�Ӽ�V�x�����i�*���S�;t�����Gt���S�\�*�`   `   ��ǽ�m����l1ջ��;��y<�j�<A�y<��;~0ջ��㼿m��ǽ#��2O����W@������1�����W@�����2O�`   `   H>%�v&ս=u���㼱@Ȼ���;,\<�\<��;�AȻ����<u��&սJ>%�^l��0����þE�⾧p���p��I�⾺�þ�0��il�`   `   Ϊ*��&ս�m��Ӽ�f�����;��$<���;8f���Ӽ�m��&սƪ*�V*|������I�����������J���ᾒ��V*|�`   `   H>%��ǽ�V�Դ�"�z�Zؚ;eך;A�z��Ӵ��V��ǽJ>%�V*|�������D����1���@���@���1�F�������O*|�`   `   $�x���^4�gm��W>�P�:S>�gm���^4�x��#�^l�������ݷ��T@�مY���b���Y��T@�ط������^l�`   `   ����N���l�n�S�0�:�N�:���S��l��N������2O��0����D���T@�#�b���v���v� �b��T@�F��ᾁ0���2O�`   `   "`̽��]���ͼ|��̄�|����ͼ��]�'`̽i�*������þI����1�مY���v�)�����v�څY���1�I����þ���i�*�`   `   ����e��{d��ם׻Ȝ׻Gd���������9I���S�W@��D�⾠����@���b���v���v���b���@����I��X@����S�=I�`   `   �T���̼_$&����M%&���̼�T�5���s�;t�����p�������@���Y� �b�څY���@�����p��
���;t��s�5��`   `   xO�ɶg�uY���X��A�g��O��ǁ�^�޽�h0����1���p�������1��T@��T@���1�����p���1�����h0�W�޽�ǁ�`   `   ����Ż5����ŻQ��7�?������'�6������I��J��F��ط�F��I��I��
������6����V���7�`   `   �
�"�����>�_^����,�9[����ｬh0�Gt�W@����þ�ᾌ�񾆭����þX@��;t��h0����*[����,��^��`   `   E7�9g�<;4H�98���#����,�X���W�޽�s���S����0������������0�������S��s�W�޽V�����,����8���`   `   +̑;�ˑ;Ĳ:����_^���6��ǁ�+5��9I�\�*��2O�il�V*|�O*|�^l��2O�i�*�=I�5���ǁ�7��^��7���.�:`   `   ��'��@�B ��bX
�q.c�u^��z�0	 ���G�f�j�1���a݅�1���q�j���G�	 �z�^��q.c�X
�C ��-A��'�`   `   �'�Ho���y������{뼭�6��F�����j��12�;���Y(��Y(�<��%2�r������F��y�6�,|�����Jy��n��(�`   `   �@��y���@���������F��:�L�t�]���3R���½yɽ�½3R��l���L�t���:�F�ɀ��������@��y��@�����`   `   C ������������������)���s�Cy��/�\=F��4S��4S�y=F��/�y��s뼘��򐙼%�����������S ���i���i��`   `   bX
��{뼧��������K��e[m���v�����ɛ�6��G��7�^ɛ������v�f[m�K������D����{�4X
�D��DJ�D��`   `   q.c���6�F�)��e[m��=��y����E����,K��J����u�E��x��=��[m����,�y�6�z.c��+���㌽�㌽�+��`   `   u^���F���:��s뼒�v��y����;XO�;�~<��<�~<XO�;��;�y����v��s���:��F���^���Dͽ!n佭��;n��Dͽ`   `   z����L�t�Cy������E�XO�; D<�o<�o<D<SP�;v�E���y�1�t����z�2��ǣ,�:M9�1M9�ã,�?��`   `   0	 �j��]����/��ɛ�����~<�o<jQ�<�o<+~<���9ɛ��/�����j�� 	 �ĤM�_�u��ሾ�፾�ሾV�u�ĤM�`   `   ��G�12�3R��\=F�7�.K���<�o<�o<@�<�J�}�y=F�&R��%2���G�~1��'}�������Dξ�Dξ����%}��w1��`   `   f�j�;���½�4S��G���J��~<D<+~<�J��G���4S��½;��p�j�τ���1ҾP����D�����D�P����1Ҿτ��`   `   1����Y(�yɽ�4S�7����VO�;RP�;���}��4S�lɽ�Y(�2���$��g���\�0G9���H���H�3G9�X�e���$��`   `   a݅��Y(��½y=F�^ɛ�x�E���;y�E�9ɛ�y=F��½�Y(�\݅��lǾg���	8�,�a��Y���	���Y��-�a��	8�e���lǾ`   `   1���<��3R���/�����x���y�����/�&R��;��2����lǾ��e G�����w�����������w�����g G����lǾ`   `   p�j�%2�l���y���v�=���v�y�����%2�p�j�$��g��e G�Ce�������߿� Xɿ�߿�����@e��e G�i��$��`   `   ��G�s��L�t��s�g[m��[m��s�1�t�j�潰�G�τ��g����	8���������<ɿ�޿�޿�<ɿ��������	8�e���Є��`   `   	 ������:����K�������:���� 	 �~1���1Ҿ\�,�a��w���߿��޿�u鿊޿�߿��w��+�a�\��1Ҿ~1��`   `   z��F��F�򐙼����,��F��z�ĤM�'}��P���0G9��Y������ Xɿ�޿�޿Xɿ�����Y��3G9�Q���%}��ȤM�`   `   �^��y�6�ɀ��&���E���y�6��^��2��_�u������D���H��	�������߿��<ɿ�߿������	����H��D�����_�u�2��`   `   q.c�,|뼶��������{�z.c��Dͽƣ,��ሾ�Dξ�����H��Y���w�����������w���Y����H�����Dξ�ሾã,��Dͽ`   `   X
�������@�����4X
��+��!n�:M9��፾�Dξ�D�3G9�-�a����@e�����+�a�3G9��D��Dξ�፾:M9�8n佫+��`   `   C ��Jy��y�S ��D���㌽���1M9��ሾ����P���X��	8�g G�e G��	8�\�Q��������ሾ:M9���콅㌽g��`   `   -A��n���@��i��DJ��㌽;n�ã,�V�u�%}���1Ҿe���e����i��e����1Ҿ%}��_�u�ã,�8n佅㌽0J��i��`   `   �'�(������i��D���+���Dͽ?��ĤM�w1��τ��$���lǾ�lǾ$��Є��~1��ȤM�2���Dͽ�+��g���i������`   `   �޻�������{���X�S���.�����-�5g�^�)��{���@ľ{����)��^#g���-�Y������S�{���؍�����`   `   ���
rH�������?9��e����½f:��'�VJ���e��9u��9u���e�VJ���'�t:���½�e��b9�C��୘��qH���`   `   ����������������U�g����ʷ���὚K����������K�����ʷ�Z����U�!���������������w��`   `   {�����）�鼿�������LB��l������~���夽�夽�~�������l��KB�*��B��U��S��C�，����_��_�`   `   X�S�?9�������L��q&�����R��>��x�#�>��$�����'��L�������_�?9�*�S��g�wn��g�`   `   ���e���U����L�缮.��PW���dx��	p���o�z�o��	p�]ex�W��M.�����*��ГU��e���������˽�˽����`   `   /�����½g���LB�q&��PW�����rMd�B�m����m�sMd����QW���&��LB�X�����½E���qF�E_#�C!)�R_#�qF�`   `   ��-�f:��ʷ��l�����dx�sMd��6`;�;��;77`;�Kd�^ex�����l��ʷ�t:���-���V�l�w�B߄�>߄�h�w���V�`   `   5g��'���Ὄ���R���	p�G�m��;G�<�;��m��	p�����������'�%g�aw�����`�ƾM:ξ`�ƾ~��aw��`   `   ^VJ��K��~��>����o�*���; �;���{�o�a���~���K�VJ�`�¾���ډ�������݉����¾`   `   �)����e�����夽x�#�{�o���m�57`;��m�{�o�[�#��夽�����e��)��V"����"?��5X��na��5X��"?����V"�`   `   {����9u����夽>���	p�wMd��Kd��	p�a���夽ۂ��9u�}���
�D>=�:�r��k�����������k��6�r�C>=�
�`   `   @ľ�9u�����~��$��^ex����_ex����~������9u�;ľ$��@�T�ۑ���@��п��ڿп�@��ۑ��>�T�$��`   `   {�����e��K��������W��QW����������K���e�|���$��6�]�����xjϿڡ��������١��zjϿ����5�]�"��`   `   �)��VJ���Ὃl�'��M.���&���l����VJ��)��
�@�T�����_�ٿ���F4&�i0�H4&����\�ٿ����C�T�
�`   `   ^��'��ʷ��KB�M�缓��LB��ʷ��'�_V"�D>=�ۑ��xjϿ���0�s`F�r`F�0����zjϿڑ��C>=�W"�`   `   #g�t:�Z���*�����*��X���t:�%g��¾��:�r��@��ڡ��F4&�s`F�\S�s`F�F4&�ڡ���@��:�r�����¾`   `   ��-���½�U�B����ГU���½��-�aw������"?��k��п���i0�r`F�s`F�j0����п�k���"?����cw��`   `   Y����e��!�V��`��e��E�����V����ډ��5X�������ڿ���H4&�0�F4&������ڿ�����5X�ډ������V�`   `   ��c9����T��?9���qF�l�w�`�ƾ����na�����п١��������ڡ��п�����na����b�ƾh�w�iF�`   `   �S�C�����C��*�S�����E_#�B߄�M:ξ����5X��k���@��zjϿ\�ٿzjϿ�@���k���5X����G:ξB߄�Q_#�����`   `   {���୘���������g��˽C!)�=߄�`�ƾ݉��"?�6�r�ۑ����������ڑ��:�r��"?�ډ�b�ƾB߄�;!)��˽�g�`   `   ؍���qH������_�wn��˽R_#�h�w�~��������C>=�>�T�5�]�C�T�C>=���������h�w�Q_#��˽cn��_�`   `   ������w���_��g�����qF���V�aw���¾V"�
�$��"��
�W"ﾡ¾cw����V�iF������g��_��w��`   `   �,W�������Ӽ�D1�r"��\�߽�%�
�h�����~�ľ��龟�r�������~�ľ����
�h��%�\�߽O"���D1�ݶӼ����`   `   ��������q演L+���������U�|�0��Ob�����E��eʦ�iʦ�F�������Ob���0��U�����í��L+��p�Ě������`   `   ��Ӽq�į���(�>S^�Ɣ�j�Ľ���aq�z�3���D��K���D�z�3�iq����]�ĽƔ�OS^���(����q漖�ӼkMμ`   `   �D1��L+���(�l�/���C�8Eg�u>���\ŽG\ܽMA�PA�V\ܽ\Ž�悔f>��pEg���C�:�/���(��L+��D1���5���5�`   `   r"�����>S^���C�iO5���4���@���T�F�i��z�����z��i���T��@���4�O5���C��S^����\"�����ja�����`   `   \�߽����Ɣ�8Eg���4�5T�
m�����j�������������Ҋ���l�T���4�pEg�Ɣ�����a�߽����Y��Y�m���`   `   �%��U�j�Ľu>����@�
m�K���������l�<*`���l�����K���
m���@�u>��[�Ľ�U��%�j�C� Y�!�`�Y�j�C�`   `   
�h�|�0����𨽀�T���������B���㻻任&������Ҋ����T��悔�����0��h�`Ǐ�2ե�f=��b=��0ե�fǏ�`   `   �����Ob�aq�\ŽF�i�j����l��㻻9ME��㻻��l�j���i�\Žsq��Ob�����"�Ⱦ�����v�������"�Ⱦ`   `   ~�ľ����z�3�G\ܽ�z�����<*`�任�㻻�)`������z�V\ܽs�3������ľL����'�{�D���U���U�~�D���'�H��`   `   ���E����D�MA齗��������l�'����l��������MA齺�D�E�����`r%���[�^���n��,����n��^����[�`r%�`   `   ��eʦ��K�PA��z������������j���z�MA��K�iʦ���b�@�.���l�����տ�m쿐m���տk���-���e�@�`   `   r��iʦ���D�V\ܽ�i�Ҋ��L���Ҋ���i�V\ܽ��D�iʦ�p���dP�U����Կ9^	�O�!��[+�O�!�9^	���ԿU���dP�`   `   ��F��z�3�\Ž��T��l�m���T�\Žs�3�E�����dP�>2��z��bn!� QL��h��h� QL�bn!�|��>2���dP�`   `   �������iq��悔�@�T���@��悔tq��������b�@�U��z��¿*���g�l��o_��l����g���*�z��U��b�@�`   `   ~�ľ�Ob����f>����4���4�u>������Ob��ľ`r%�.�����Կbn!���g��Q������ߝ���Q����g�bn!���Կ-���ar%�`   `   ������0�]�ĽpEg�O5�pEg�[�Ľ��0�����L����[�l���9^	� QL�l��������������l�� QL�9^	�l�����[�L��`   `   
�h��U�Ɣ���C���C�Ɣ��U��h�"�Ⱦ��'�^����տO�!��h�o_��ߝ������p_���h�O�!���տ^����'�$�Ⱦ`   `   �%�����OS^�:�/��S^������%�`Ǐ����{�D��n���m��[+��h�l���Q��l���h��[+��m��n��{�D����`Ǐ�`   `   \�߽í���(���(����a�߽j�C�2ե�����U�,����m�O�!� QL���g���g� QL�O�!��m�,�����U���0ե�b�C�`   `   O"���L+�����L+�\"����� Y�f=��v����U��n����տ9^	�bn!���*�bn!�9^	���տ�n����U�s��f=��Y����`   `   �D1��p�q漣D1�����Y�!�`�b=����~�D�^��k�����Կ|��z�꿷�Կl���^��{�D���f=���`��Y���`   `   ݶӼĚ����Ӽ��5�ja���Y�Y�0ե���񾐸'���[�-���U��>2��U��-�����[���'����0ե�Y��Y�`a����5�`   `   ��������kMμ��5����m���j�C�fǏ�"�ȾH��`r%�e�@��dP��dP�b�@�ar%�L��$�Ⱦ`Ǐ�b�C��������5�6Mμ`   `   k��������!�Z^a�c��V�*[N�G���zľ�5��y���T'��-��T'�|���5��zľG���<[N�V��b��[^a��!�����`   `   ����$$ݼ�N�?\��	���뽼,%�t�^�n���ȭ�#�ƾ�Ծ�Ծ$�ƾ�ȭ�o����^��,%����	��_\��N�$ݼ���`   `   �!��N��N0�=�[�͏��k���D���T!��E�[�e��|�����|�[�e��E��T!��D���k��"͏�=�[��N0��N��!���`   `   [^a�?\�=�[�ȣg��@��|I���Ժ��\�������������������\ཚԺ��I���@����g�#�[�_\�d^a���e���e�`   `   c���	��͏��@����x�Ģ~����dt������E����ζ�E�������dt��:���Ģ~�o�x��@��?͏��	���b��������ƽ����`   `   V����k��|I��Ģ~�4�^�Q��8P�'�T���X���X�4�T��8P��Q��^��~��I���k����V��(�V6'�S6'��(�`   `   *[N��,%��D���Ժ����Q�nj)�e������	����e��mj)�Q�����Ժ��D���,%�3[N��os�f����i��k����os�`   `   G���t�^��T!��\�dt���8P�e����#
˼>
˼	��J���8P�tt���\��T!���^�H����)���о+�߾'�߾�о�)��`   `   zľn���E��������'�T����#
˼޳��#
˼܎�'�T�}������%�E�n��zľrD�����-� 4��-���rD��`   `   �5���ȭ�[�e���E�����X��	�>
˼$
˼�	���X�U������T�e��ȭ��5���3*���X�(s��j��k��*s����X��3*�`   `   y��#�ƾ�|�����ζ���X����	��܎���X��ζ�����|�#�ƾ{��!{V�2���L�����ѿ)ܿ��ѿL���4���!{V�`   `   �T'��Ծ������E���4�T�e��J��'�T�U����������Ծ�T'�|�Q/��S^�d��n&�o&�e��Q^�P/��|�`   `   �-��Ծ�|���������8P�mj)��8P�}�������|��Ծ߿-������Ͽ(L�*�E���n��|���n�+�E�(L��Ͽ����`   `   �T'�$�ƾ[�e����dt���Q�Q�tt�����T�e�#�ƾ�T'�����}2ٿ�h%��Yn��;��+͹�*͹��;���Yn��h%�}2ٿ����`   `   |���ȭ��E��\�:����^�����\�%�E��ȭ�{��|��Ͽ�h%�b�~�<����l���5��l��<���a�~��h%��Ͽ|�`   `   �5��o���T!��Ժ�Ģ~��~��Ժ��T!�n���5��!{V�Q/��(L��Yn�<���-�*u$�*u$�-�<����Yn�(L�P/��"{V�`   `   zľ��^��D���I��o�x��I���D����^�zľ�3*�2���S^�*�E��;���l��*u$���6�*u$��l���;��*�E�S^�2����3*�`   `   G����,%��k���@���@���k���,%�H���rD����X�L���d����n�+͹��5�*u$�*u$��5�*͹���n�e��L�����X�tD��`   `   <[N���"͏���g�?͏���3[N��)����(s����ѿn&��|�*͹��l��-��l��*͹��|�n&���ѿ(s�����)��`   `   V��	��=�[�$�[��	��V��os��о�-�j��)ܿo&���n��;��<���<����;����n�n&�)ܿk���-��о�os�`   `   �b��_\��N0�_\��b���(�f���+�߾ 4�k����ѿe��+�E��Yn�a�~��Yn�*�E�e����ѿk�� 4�+�߾k����(�`   `   [^a��N��N�d^a�����V6'��i��'�߾�-�*s��L���Q^�(L��h%��h%�(L�S^�L���(s���-�+�߾�i��S6'�����`   `   �!�$ݼ�!���e���ƽS6'�k����о����X�4���P/���Ͽ}2ٿ�ϿP/��2�����X����оk���S6'���ƽ��e�`   `   �����������e������(��os��)��rD���3*�!{V�|���������|�"{V��3*�tD���)���os��(�������e�ȓ�`   `   �����ༀ�&��τ�,ӽQ�"�;�q�,����V�;���3���H�Y�P���H��3�;���V�,���J�q�Q�"�ӽ�τ���&����`   `   ����w��D6�Fk������:�$�C��������Ͼ0��:���:��0��Ͼ�������C��:�����Sk���D6��w���`   `   ��&��D6���U�����z���Z�轠���DC�p�n��ኾ.b��&<��*b���ኾw�n��DC����Z�����������U��D6��&���!�`   `   �τ�Fk�������w�����^ý�[�8����$�x 7�bMA�dMA�~ 7���$�.���[�tý���~w������Sk���τ�M���R���`   `   ,ӽ���z������T���vʩ�Tm����Ͻ�D�r9����r9�D住�Ͻsm��vʩ�1�������������ӽ���Q潊�`   `   Q�"��:�Z��^ývʩ��>������/��0*��s9��o9��5*���/������>���ʩ�týN���:�T�"�M6��cA��cA��L6�`   `   ;�q�$�C�����[�Tm�����S��~8��b��b�`��~8��S�����Ym���[콛��$�C�B�q��ƍ�����  �������ƍ�`   `   ,�������DC�8����Ͻ�/��~8����i�r^�r^���i�s8���/����Ͻ.���DC����.���Z\Ӿn$��Oj�Nj�m$��_\Ӿ`   `   �V����p�n���$��D�0*��b��r^���S�r^�q��0*���D位�$���n�����V辩~���6�N�	�V�N���6��~�`   `   ;���Ͼ�ኾx 7�r9�s9��b�r^�r^�V�o9���9�~ 7��ኾ�Ͼ;��[sK�v���C����c���c��D���v���YsK�`   `   �3�0�.b��bMA����o9��a����i�r��o9��׮��bMA�.b��0�3�Od��ޟ���k�����	����k�ߟ��Od��`   `   ��H��:��&<��dMA�r9�5*��8��s8��0*���9�bMA�$<���:����H�[8��[�޿uS�8y?�\qX�]qX�8y?�tS�[�޿\8��`   `   Y�P��:��*b��~ 7��D��/��S���/���D�~ 7�.b���:��W�P�3>���Y���>��M���}��Y	���}���M����>��Y�3>��`   `   ��H�0��ኾ��$���Ͻ��������Ͻ��$��ኾ0��H�3>���(�S:W�D-��������������D-��S:W��(�2>��`   `   �3��Ͼw�n�.��sm���>��Ym��.����n��Ͼ�3�[8���Y�S:W�P����q�>��OS�>��q�P���S:W��Y�[8��`   `   ;������DC��[�vʩ��ʩ��[��DC����;��Od��[�޿��>�D-���q�RES���������RES��q�D-����>�[�޿Od��`   `   �V�������tý1���tý�������V�[sK�ޟ��uS��M������>������M������>������M��uS�ޟ��[sK�`   `   ,����C�Z��������O��$�C�.����~�v����k�8y?��}�����OS����������OS����}��8y?��k�v����~�`   `   J�q��:�����~w�������:�B�q�Z\Ӿ��6�C�����\qX�Y	����>�RES�>���Z	��\qX���C�����6�Z\Ӿ`   `   Q�"����������������T�"��ƍ�n$��N��c����	�]qX��}�������q��q������}��\qX���	��c��N�m$���ƍ�`   `   ӽSk����U�Sk��ӽM6�����Oj�	�V��c����8y?��M��D-��P���D-���M��8y?����c���V�Oj�����M6�`   `   �τ��D6��D6��τ��ὠcA�����Nj�N�D����k�tS���>�S:W�S:W���>�uS��k�C���N�Oj������cA���`   `   ��&��w��&�M����Q潞cA�����m$����6�v���ߟ��[�޿�Y��(��Y�[�޿ޟ��v�����6�m$�������cA��Q�M���`   `   �������!�R������L6��ƍ�_\Ӿ�~�YsK�Od��\8��3>��2>��[8��Od��[sK��~�Z\Ӿ�ƍ�M6���M�����!�`   `   KEڼ����,;�1ړ�W��0�3�e��ʽ��� �7^%��|G��,`��>i��,`��|G�7^%��� �ʽ�e��0�3�B��1ړ�$,;�����`   `   ������]O�r-��j�ٽ�	��\��V��ʾ��e��%�o��p���%��e�ʾ��V���\��	�u�ٽ|-���]O������`   `   ,;��]O�тv�>���/z̽���1�B_b�������3s��Q���/s��������B_b��1���3z̽>���тv��]O�,;��5�`   `   1ړ�r-��>����]����ƽ`^�
=�7�-���H�=�^���j���j�B�^���H�/�-�=�q^ｒ�ƽ�]��4���|-��6ړ�>=��@=��`   `   W��j�ٽ/z̽��ƽ��̽�kݽ�)��Wz
��W�Y)"���%�Y)"��W�Wz
��)���kݽĆ̽��ƽHz̽j�ٽI���O������O��`   `   0�3��	���`^��kݽ�\ٽm�߽,��{���������~���7��d�߽x\ٽ�kݽq^����	�2�3��G�=R�=R��G�`   `   e���\��1�
=��)��m�߽�v׽~׽�*ڽK�۽�*ڽ~׽�v׽m�߽�)��
=��1��\�e��m������!J������m��`   `   ʽ��V��B_b�7�-�Wz
�,��~׽VϽ��̽��̽VϽ~׽7��]z
�/�-�=_b��V�� ʽ�"���	������&�`   `   �� �ʾ������H��W�{����*ڽ��̽�[ɽ��̽�*ڽ{����W���H����ʾ��� �i&���I��{c�m��{c��I�i&�`   `   7^%��e����=�^�Y)"����K�۽��̽��̽C�۽���_)"�B�^�����e�8^%�$�a�E��ߩ��������ߩ��E��!�a�`   `   �|G��%�3s����j���%�����*ڽVϽ�*ڽ�����%���j�3s���%��|G��]��8<ƿ����X��~��W������9<ƿ�]��`   `   �,`�o��Q�����j�Y)"����~׽~׽{���_)"���j�N���p���,`�3���]���.�<^�M}�M}�<^��.�]��4���`   `   �>i�p��/s��B�^��W�8�뽲v׽8���W�B�^�3s��p���>i�컿�R���]�)P���]�������]��)P����]��R�컿`   `   �,`��%������H�Xz
�d�߽m�߽]z
���H�����%��,`�컿�p��|����$T��2��2�#T�����|��p�컿`   `   �|G��e辷��/�-��)��x\ٽ�)��/�-�����e��|G�3����R��|�!����}2��7u��Z���7u��}2�!����|��R�3���`   `   7^%�ʾ�B_b�=��kݽ�kݽ=�=_b�ʾ�8^%��]��]����]�����}2�<U���u���u��<U���}2������]�]���]��`   `   �� ��V���1�r^�Ć̽r^��1��V���� �$�a�8<ƿ�.�)P��$T��7u��u��[���u���7u�$T�)P���.�8<ƿ$�a�`   `   ʽ��\�����ƽ��ƽ���\� ʽ�i&�E������<^��]���2��Z���u���u���Z���2��]��<^�����E��j&�`   `   e���	�4z̽�]��Hz̽�	�e��"辁�I�ߩ��X��M}������2��7u�<U���7u��2�����M}�W��ߩ����I�"�`   `   0�3�v�ٽ>���4���k�ٽ2�3�m�����{c����~��M}��]��#T��}2��}2�$T��]��M}�~������{c���k��`   `   B��|-��҂v�|-��I�齟G�����	��m����W��<^�)P�����!������)P��<^�W�����m�	�������G�`   `   1ړ��]O��]O�6ړ��O��=R�!J�����{c�ߩ�������.���]��|��|���]��.�����ߩ���{c�	��J��=R��O��`   `   $,;��,;�>=�����=R��������I�E��9<ƿ]���R��p��R�]��8<ƿE����I�������=R����>=��`   `   ���������5�@=���O���G�m��&�i&�!�a��]��4���컿컿3����]��$�a�j&�"�k���G��O��>=���5�`   `   ���`gJ��=�����K�=�����tfƾ#2��,�uBO�K�h�mr�K�h�vBO��,�"2�tfƾ����K�=�����=��ngJ����`   `   ����(��ud�^<����+�� n�~����̾�������"��#����������̾����� n��
+���d<���ud��(����`   `   `gJ��ud�������Zq��I��YJ�����ᚾ���0þFɾ�0þ���ᚾ����YJ��I�]q��������ud�YgJ��KB�`   `   �=��^<������"ʽF ����H1��!S��&s�.���$���$��.���&s��!S��H1���M �"ʽ���d<���=��[G��\G��`   `   �����Zq�F �8�xz��$��9���K�غX��\]�غX���K��9��$�xz��7�F �kq�������] ���] �`   `   K�=�+��I���xz��H��
!�D~-��38�'Y>�$Y>��38�I~-��
!��H�{z����I��
+�M�=�%2N���W���W�"2N�`   `   ����� n��YJ��H1��$��
!���$��1+��0���2��0��1+���$��
!��$��H1��YJ�� n������������9����������`   `   tfƾ~�������!S��9�D~-��1+�n-���.���.�l-��1+�I~-��9��!S��������ufƾ���}�����ߖ�}�����`   `   #2��̾�ᚾ�&s���K��38��0���.�1�.���.��0��38���K��&s��ᚾ�̾!2��*�N��h�ïq��h�N��*�`   `   �,�������.��غX�'Y>���2���.���.���2�%Y>�ܺX�.��볲������,��5h�*���Y���~�¿~�¿Z���*����5h�`   `   uBO�����0þ�$���\]�%Y>��0�l-��0�%Y>��\]��$���0þ���vBO�ނ���:˿T��-B��� �-B�T���:˿ނ��`   `   K�h�"��Fɾ�$��غX��38��1+��1+��38�ܺX��$��Dɾ#��K�h�R���ۈ��^3�ܵd�Ԇ��Ԇ��ܵd��^3�ۈ�S���`   `   mr�#���0þ.����K�I~-���$�I~-���K�.���0þ#��kr�d��Hd��d�����)������)�������d�Hd�d��`   `   K�h�������&s��9��
!��
!��9��&s�볲����K�h�d��q��~��b�������:��:����b�����q��d��`   `   vBO������ᚾ�!S��$��H��$��!S��ᚾ����vBO�R���Hd�~���p����:�.M������.M����:��p��~��Hd�R���`   `   �,��̾����H1�xz�|z��H1�����̾�,�ނ��ۈ��d�b�����:������5���5��������:�b����d�ۈ�߂��`   `   "2������YJ����7����YJ�����!2��5h��:˿�^3��������.M���5��U���5��.M����������^3��:˿�5h�`   `   tfƾ� n��I�N �G ��I�� n�ufƾ�*�*���T��ܵd�)���:������5���5�������:�)��ܵd�T��*����*�`   `   �����
+�]q꽍"ʽkq��
+��������N�Y���-B�Ԇ�������:�.M������.M���:�����Ԇ��-B�Y���N����`   `   K�=�����������M�=����}���h�~�¿�� �Ԇ��)�������:���:����)��Ԇ���� �~�¿�h�}�����`   `   ���d<�����d<�����%2N��������ïq�~�¿-B�ܵd�����b����p��b�������ܵd�-B�~�¿ïq��������%2N�`   `   �=���ud��ud��=���] ���W�9���ߖ��h�Z���T���^3��d���~���d��^3�T��Y����h����7�����W��] �`   `   ogJ��(�YgJ�[G�����W�����}��N�*����:˿ۈ�Hd�q��Hd�ۈ��:˿*���N�}��������W��[G��`   `   �������KB�\G���] �"2N��������*��5h�ނ��S���d��d��S���߂���5h��*�������%2N��] �[G���KB�`   `   �a�`��Q-X��C���q ���A�yq���bƾ���'%)��J�5�b�qk�5�b��J�'%)�����bƾzq����A��q ��C��T-X�`��`   `   `��Ii7��,z�Cp��Cm�'u7�Fa|�L����Ӿc�����{x�|x���a�����ӾM��Fa|�&u7�Dm�Dp���,z�Ki7�e��`   `   Q-X��,z�lڛ��8˽�����1��e�8������� �ži�־D�ܾe�־ �ž����8����e���1�����8˽nڛ��,z�I-X��^M�`   `   �C��Cp���8˽���>��mZ4��n[�{+��5��uʣ�0׫�1׫�wʣ�5��y+���n[�pZ4�?�����8˽Dp���C��;���:���`   `   �q �Cm����>����%�Ж?��b]��y{����>���I���>�������y{��b]�Ж?���%�?�����Cm��q �I�\��I�`   `   ��A�'u7���1�mZ4�Ж?�TDR�'i���� "��h8��g8�� "�����'i�PDR�і?�pZ4���1�&u7���A�V�L��S��S�U�L�`   `   yq��Ea|��e��n[��b]�'i��2z��B拾�+��D拾��2z�'i��b]��n[��e�Fa|�yq�����X慨�T��X慨���`   `   �bƾL��8���{+���y{���������p:��o:�����������y{�y+��7���M���bƾ��较����������`   `   �����Ӿ����5����� "��B拾p:��Ơ��p:��D拾 "�����5��������Ӿ���|�$�lD��;[���c��;[�kD�|�$�`   `   '%)�c��� �žuʣ�>���h8���+��o:��p:���+��g8��?���wʣ��ža���'%)��^��u���N��7���7����N���u���^�`   `   �J���h�־0׫�I���g8��D拾����D拾g8��J���0׫�g�־��	�J�Yo��B���}U����)���}U�B���Yo��`   `   5�b�{x�D�ܾ1׫�?��� "���� "��?���0׫�C�ܾ|x�5�b��~���[��$�WP���k���k�WP���$��[��~��`   `   qk�|x�e�־wʣ��������2z�������wʣ�h�־|x�qk��۶�=`�h�O�-r��yȵ����yȵ�-r��h�O�<`��۶�`   `   5�b��� �ž5���y{�'i�'i��y{�5���ž��5�b��۶�����mk�����=�z/�z/��=�����mk�����۶�`   `   �J�a�������y+���b]�PDR��b]�y+������a���	�J��~��=`��mk��|��P���Y��?r���Y�P��|���mk�=`��~��`   `   '%)���Ӿ8����n[�Ж?�і?��n[�8�����Ӿ'%)�Yo���[�h�O����P�)8r���������)8r�P����h�O��[�Yo��`   `   ���M���e�pZ4���%�pZ4��e�M������^�B�����$�-r���=���Y�����c[��������Y��=�-r����$�A����^�`   `   �bƾFa|���1�@��?����1�Fa|��bƾ|�$��u��}U�WP�yȵ�z/��?r����������?r�z/�yȵ�WP�}U��u��{�$�`   `   zq��&u7���������&u7�yq�����lD��N������k����z/���Y�)8r���Y�z/������k����N��lD����`   `   ��A�Dm��8˽�8˽Cm���A�������;[�7����)���k�yȵ��=�P�P��=�yȵ���k��)�7����;[������`   `   �q �Dp��nڛ�Dp���q �V�L�X慨����c�7�����WP�-r������|�����-r��WP���7�����c���W慨V�L�`   `   �C���,z��,z��C��I��S��T�����;[��N��}U��$�h�O��mk��mk�h�O���$�}U�N���;[����T���S�I�`   `   U-X�Ki7�J-X�;���\���S�X慨��kD��u��B����[�<`����=`��[�A����u��lD���W慨�S�[��;���`   `   `��f���^M�:���I�U�L�������|�$��^�Yo���~���۶��۶��~��Yo���^�{�$���辋��V�L�I�;����^M�`   `   ����(�vJj�뿯�g���TD�P���ͯ��c���Z ��>��&S���Z��&S��>�Z �e���ͯ��N����TD�j��뿯�nJj��(�`   `   �(��wL�1����'ǽ�FmF��E��+���0cھ���6��^��^��6���.cھ+����E��GmF���'ǽ3����wL��(�`   `   vJj�1������Q�����wP��v�����Oľj�޾��[�����j�޾Rľ����v���wP����Q����1���pJj�Y�[�`   `   뿯��'ǽQ�����.�7���d������Y��������ξ�Qؾ�Qؾ��ξ�����Y��������d�+�7����S��'ǽ쿯��ऽ�ऽ`   `   f�����.�7���Y�ٹ���n��Γ���F����;b8Ҿ��;�F��Γ���n��ٹ����Y�.�7����h��q ��{��q �`   `   �TD�FmF��wP���d�ٹ�������?�����̾�*վ�*վ��̾@����󩾙��ع����d��wP�GmF��TD��ZF���H���H��ZF�`   `   P����E���v�������n����A��,ξN�پ�0޾Q�پ,ξ>���󩾽n�������v���E��P���!3��=~���S��<~��!3��`   `   ͯ��+�������Y��Γ��?���,ξܾF��E��
ܾ,ξ@���͓���Y�����+���ί���ؾR?�������S?��ؾ`   `   c���0cھOľ�����F����̾N�پF��̴�F��N�پ��̾�F������Oľ0cھc����g�X/�oeA��#H�oeA�X/��g�`   `   Z ���j�޾��ξ��;�*վ�0޾E��F�㾿0޾�*վ��;��ξk�޾��Z ��fI�iJw���uG��uG����iJw��fI�`   `   �>��6���Qؾb8Ҿ�*վQ�پ
ܾN�پ�*վe8Ҿ�Qؾ��6��>�P�|��A��)ͿJ쿹���K�)Ϳ�A��P�|�`   `   �&S��^�[����Qؾ��;��̾,ξ,ξ��̾��;�Qؾ[����^��&S�0`����ο��	��*���>���>��*���	���ο0`��`   `   ��Z��^��𾷗ξ�F��@���>��@����F����ξ��^���Z��+���:*���d�ݖ��1��ݖ����d��:*����+��`   `   �&S��6�j�޾����Γ���󩾆�͓������k�޾�6��&S��+�����`�>�����q��O���O���q������`�>�����+��`   `   �>���Rľ�Y���n������n���Y��Oľ���>�0`����`�>����������"��q'��"���������`�>���0`��`   `   Z �.cھ�������ٹ��ع���������0cھZ �P�|���ο�:*���������cm'��lN��lN�cm'����������:*���οQ�|�`   `   e���+����v����d���Y���d��v��+���c����fI��A����	���d�q���"��lN��xe��lN��"�q����d���	��A���fI�`   `   ͯ���E���wP�,�7�.�7��wP��E��ί���g�iJw�)Ϳ�*�ݖ��O����q'��lN��lN��q'�O���ݖ���*�)ͿiJw��g�`   `   N���GmF���������GmF�P����ؾX/���J���>�1��O����"�cm'��"�O���1����>�J���X/��ؾ`   `   �TD��Q��S����TD�!3��R?�oeA�uG��������>�ݖ��q����������q��ݖ����>�����uG��neA�S?�#3��`   `   j���'ǽ����'ǽh���ZF�=~������#H�uG��K��*���d���������������d��*�J�uG���#H����;~���ZF�`   `   뿯�3���1���쿯�q ���H��S�����oeA���)Ϳ��	��:*�`�>�`�>��:*���	�)Ϳ��neA�����S����H�q �`   `   nJj��wL�qJj��ऽ�{����H�<~��S?�X/�iJw��A����ο�������ο�A��iJw�X/�S?�;~����H��{���ऽ`   `   �(��(�Z�[��ऽq ��ZF�!3���ؾ�g��fI�P�|�0`���+���+��0`��Q�|��fI��g��ؾ#3���ZF�q ��ऽ^�[�`   `   oM-��<C�Z����(���V��)J��3��3(��Ƨ���\���0�H�B��#I�H�B���0��\�˧��3(���3���)J��V��(��O����<C�`   `   �<C��l�A��cM��� ��+]�����h��h�ɳ�B[�X  �X  �C[�ɳ��g��h������+]��� �]M�A���l��<C�`   `   Y���A��&Խ�l��{@�_�|������*žnD�z��p���Z�o��z��qD��*ž����_�|��{@��l�%ԽA��Y���%�s�`   `   �(��cM��l�78��^l�������-پ����ʈ�������ˈ������-پ������^l�78��l�\M佡(��eN��bN��`   `   �V��� ��{@��^l�`������`$վ(^���
	��>��x��>��
	�(^��]$վ����d���^l��{@��� ��V����0����`   `   �)J��+]�_�|����������Ծ� �����X��������X���� ����Ծ�������c�|��+]��)J��m@�Q�<�S�<��m@�`   `   �3�����������`$վ� ��{�g[�M&��)�M&�g[�}{�� ��c$վ����������3���|��Xэ����Vэ��|��`   `   3(���h���*ž�-پ(^����g[��)��/��/��)�i[���%^���-پ�*ž�h��2(��;�ƾ&�Ѿr�ؾs�ؾ'�Ѿ9�ƾ`   `   Ƨ��h�nD������
	��X�M&��/��Y3��/�M&��X��
	�����lD�h�ȧ��K��dN���!��a&���!�eN�K��`   `   �\�ɳ�z��ʈ��>�����)��/��/��)�����>�ˈ�{��ɳ��\�V�0��O���j�Ș{�Ș{���j��O�V�0�`   `   ��0�B[�p������x����M&��)�M&�����x����o��B[���0�
�Y�xi��eآ�_�����`��eآ�wi��
�Y�`   `   H�B�X  ��Z�����>��X�g[�i[��X��>�����Z�X  �G�B��e|��6��B�ԿW ��{��{�W �B�Կ�6���e|�`   `   �#I�X  �o��ˈ��
	���}{����
	�ˈ�o��X  ��#I�`���&��� �s&�E��#Q�E�s&�� ��&��`��`   `   H�B�C[�z������(^��� ��� ��&^������{��B[�G�B�`��=�ſ���`qE��}��������}�_qE����>�ſ`��`   `   ��0�ɳ�qD辮-پ]$վ��Ծc$վ�-پlD�ɳ���0��e|��&������Q��(��`��@M��`���(���Q�����&���e|�`   `   �\��g��*ž�������������*žh��\�
�Y��6��� �`qE��(���N��+_��+_���N���(��_qE�� ��6���Y�`   `   ˧���h���������e����������h��ȧ��V�0�xi��B�Կs&��}�`��+_��7��+_��`���}�s&�B�Կwi��V�0�`   `   3(�����`�|��^l��^l�d�|����2(��K���O�eآ�W �E����@M��+_��+_��@M�����E�W �eآ��O�J��`   `   �3���+]��{@�78��{@��+]��3��;�ƾdN���j�_���{��#Q����`���N��`������#Q��{�_����j�eN�;�ƾ`   `   �)J��� ��l��l��� ��)J��|��&�Ѿ��!�Ș{�����{�E��}��(���(���}�E��{����Ș{���!�'�Ѿ�|��`   `   �V�]M�&Խ]M��V��m@�Xэ�r�ؾ�a&�Ș{�`��W �s&�_qE��Q�_qE�s&�W �_��Ș{��a&�r�ؾTэ��m@�`   `   �(��A��A���(����Q�<����s�ؾ��!���j�eآ�B�Կ� �������� �B�Կeآ���j���!�r�ؾ���S�<���`   `   O����l�Y���fN���0��S�<�Vэ�'�ѾeN��O�wi���6���&��>�ſ�&���6��wi���O�eN�'�ѾTэ�S�<��0��fN��`   `   �<C��<C�%�s�bN�����m@��|��9�ƾK��V�0�
�Y��e|�`��`���e|��Y�V�0�J��;�ƾ�|���m@���eN��5�s�`   `   �S��&k������Vؽ�;��MX�'P��_����������7*� �9�U?� �9��7*�������_���P���MX��;��Vؽ�����&k�`   `   �&k��Z��D���Ɇ�#�<�YO���g����ԾA�����%��\.��\.���%�	��?���Ծ�g��]O���<�Ć�R����Z���&k�`   `   ����D���n���1��Mp���E�Ⱦԓ��m,���!�+�-��2�)�-���!�o,�ԓ��C�Ⱦ���Mp��1�l��D��������ƌ�`   `   �VؽɆ��1��k�4���V�ž����b��4�&�#�6�s�>�u�>�$�6�2�&�b������S�ž/����k��1�Ć��Vؽj���g���`   `   �;�#�<��Mp�4���vrž�����S���-� �A���N��gS���N�"�A���-��S�����~rž4����Mp�#�<��;��k�� ��k�`   `   �MX�YO����V�ž�������rj2�w�J�_�\���e���e�]�\�x�J�tj2��������S�ž��]O���MX��@��4��4��@�`   `   'P���g��E�Ⱦ�����S�rj2�U�M��6d��r�d�w�"�r��6d�R�M�rj2��S�����E�Ⱦ�g��%P��?��{��ȹ�x��?��`   `   _�����Ծԓ��b����-�w�J��6d��Hw�� ��Hw��6d�x�J���-�b��ؓ����Ծ^����x��1ȷ��K���K��2ȷ��x��`   `   ���A�m,�4�&� �A�_�\��r���[����r�_�\�"�A�4�&�k,�A�����������B!���������`   `   �������!�#�6���N���e�d�w� ��f�w���e���N�$�6���!�	�����q���*�l�8�,"B�+"B�k�8��*�r��`   `   �7*���%�+�-�s�>��gS���e�"�r��Hw��r���e��gS�s�>�(�-���%��7*�wD<�ƣX��.x����PU������.x�ģX�wD<�`   `    �9��\.��2�u�>���N�]�\��6d��6d�_�\���N�s�>��2��\.���9�^�V�."�������E����ƿ��ƿ�E������."��]�V�`   `   U?��\.�)�-�$�6�"�A�x�J�R�M�x�J�"�A�$�6�(�-��\.�U?���e������຿�e�Ol�c�Ol��e��຿������e�`   `    �9���%���!�2�&���-�tj2�rj2���-�4�&���!���%���9���e�)՗�0̿\��-#��5��5��-#�\�0̿*՗���e�`   `   �7*�	��o,�b���S�����S�b��k,�	���7*�^�V�����0̿�E��[6�|7Y��g�{7Y��[6��E�0̿����^�V�`   `   ���?�ԓ������������������ؓ��A����wD<�."���຿\��[6��.g����������.g��[6�\��຿."��yD<�`   `   �����ԾC�ȾS�ž~ržS�žE�Ⱦ��Ծ���q��ƣX������e濩-#�|7Y�����A�������|7Y��-#��e濅���ģX�q��`   `   `����g����/���4����򝾥g��^�������*��.x��E��Ol��5��g����������g��5�Ol��E���.x��*����`   `   P��]O���Mp��k��Mp�]O��%P���x�����l�8������ƿc��5�{7Y��.g�|7Y��5�b���ƿ���l�8������x��`   `   �MX��<��1��1�#�<��MX�?��1ȷ��,"B�PU����ƿOl��-#��[6��[6��-#�Ol���ƿQU��+"B��2ȷ�?��`   `   �;�ņ�l��ņ��;��@�{���K��B!�+"B�����E���e�\��E�\��e濺E�����+"B�E!��K��u���@�`   `   �VؽS���D����Vؽ�k��4�ȹ��K���k�8��.x������຿0̿0̿�຿�����.x�l�8���K��ӹ��4��k�`   `   �����Z������k���� ��4�x��2ȷ������*�ģX�."������*՗�����."��ģX��*�����2ȷ�u���4�� �k���`   `   �&k��&k��ƌ�g����k��@�?���x�����r��wD<�]�V���e���e�^�V�yD<�q������x��?���@��k�j����ƌ�`   `   xǃ��ܐ��˸��\��Z0�nr�����ߔо���;�P/��=�(�B��=�P/�;����ߔо����nr�0Z0��\���˸��ܐ�`   `   �ܐ�8䮽�����$�cEd�������Ⱦ�(��<���=/�Z�@���J���J�\�@��=/�9���(���Ⱦ����UEd���$���:䮽�ܐ�`   `   �˸�����o!��|_����G ɾ. ���yW8�۫N�(J]�t_b�&J]�۫N�{W8���. �G ɾ����|_��o!�����˸�;�`   `   �\����$��|_��旾1�ʾW�9�#���C���_��6t����6t���_���C�<�#�W�*�ʾ�旾�|_���$��\���ؽ�ؽ`   `   Z0�cEd����1�ʾU���i(��
M��zn�u���R���`���R���v����zn��
M��i(�[��1�ʾ���cEd�&Z0��V�6���V�`   `   nr�����G ɾW��i(��gP�S�v��&��y���x(��w(��w����&��W�v��gP��i(�W�M ɾ����ir���H��>5��>5���H�`   `   ������Ⱦ. �9�#��
M�S�v��ڎ������r��կ��r�������ڎ�S�v��
M�9�#�. ���Ⱦ����&����u��'m��u�&���`   `   ߔо�(������C��zn��&������ͥ��I��G��̥�������&���zn���C���(��ܔоVU���o��� ��� ���o��RU��`   `   ���<��yW8���_�u���y����r��I���6��I���r��y���v�����_�uW8�<�����G�{{ݾj�پR�ؾj�پ{ݾG�`   `   ;��=/�۫N��6t�R���x(��կ�G��I��կ�w(��Q����6t�ޫN��=/��:�EN�������X��X������FN�`   `   P/�Z�@�(J]��`���w(���r��̥���r��w(��c����%J]�Z�@�P/��*�a�0�na<�D9G� �K�H9G�na<�_�0��*�`   `   �=���J�t_b��R���w�����������y���Q����w_b���J��=��u?� [O��h����]b��\b�����h� [O��u?�`   `   (�B���J�&J]��6t�v����&���ڎ��&��v����6t�%J]���J�)�B��K��'e�z��P������:д����P���z���'e��K�`   `   �=�\�@�۫N���_��zn�W�v�S�v��zn���_�ޫN�Z�@��=��K��m�d%��{c����Ͽ���⿝�Ͽzc��d%���m��K�`   `   P/��=/�{W8���C��
M��gP��
M���C�uW8��=/�P/��u?��'e�d%���'��"�㿤���	����"���'��d%���'e��u?�`   `   ;�9����<�#��i(��i(�9�#���<���:��*� [O�z��{c��"�㿩J	��������J	�!��zc��z�� [O��*�`   `   ����(��. �W�[��W�. ��(�����EN�a�0��h�P�����Ͽ������' ���������ϿQ����h�_�0�EN�`   `   ߔо�ȾH ɾ*�ʾ1�ʾM ɾ��ȾݔоG����na<����������	��������	���������pa<����G�`   `   ������������旾�����������WU��{{ݾ��E9G�]b��:д��⿣���J	������9д�]b��D9G����{ݾWU��`   `   nr�UEd��|_��|_�dEd�ir�&����o��j�پ�X� �K�\b�������Ͽ"��!�㿜�Ͽ���]b��"�K��X�d�پ�o��.���`   `   0Z0���$��o!���$�&Z0���H��u�� ��R�ؾ�X�H9G����P���zc���'��zc��Q������D9G��X�[�ؾ� ���u���H�`   `   �\��������\���V��>5��'m�� ��j�پ��na<�h�z��d%��d%��z���h�pa<���d�پ� ���'m��>5��V�`   `   �˸�;䮽�˸��ؽ6���>5��u��o��{ݾ���_�0� [O��'e��m��'e� [O�_�0�����{ݾ�o���u��>5�C���ؽ`   `   �ܐ��ܐ�;��ؽ�V���H�&���RU��G�GN��*��u?��K��K��u?��*�EN�G�WU��.�����H��V��ؽP�`   `   T���ҝ���ང���N���a����e�Y|�h�+���A�8�P�ۯU�8�P���A�h�+�`|��e�R�����"�N������ҝ��`   `   ҝ��q׽����qI�WN��޻�J������8��eT�f�h���s���s�i�h��eT��8����T��޻�MN���qI����r׽ĝ��`   `   �འ���H�ҋ��쿾א���#�3�H�n�j��6��9���a��
9���6��q�j�3�H�	�#�א���쿾ҋ��H�������ʽ`   `   ����qI�ҋ����,�R�+���V����ȑ������������������ȑ���ƇV�P�+�,����ҋ��qI�|���N���N��`   `   �N�WN���쿾,�sr.��F^�����͝��d�������[ǿ�����d���͝�����F^�zr.�,��쿾WN���N�C<%�6��C<%�`   `   ��޻�֐��R�+��F^�ϡ��>¤�|�����ٿ�?��?鿎�ٿ|���A¤�С���F^�P�+�ސ��޻�
����[��?��?���[�`   `   a���J���#���V����>¤���ſگ�nW����pW�گ迼�ſ>¤������V�
�#�J��_���x����v��kh���v�x��`   `   �e쾼��3�H����͝�|���گ���'��&����ݯ�|����͝���7�H�����e�邼��柾A���E����柾䂼�`   `   Y|��8�n�j��ȑ��d����ٿnW�'��J��'��nW���ٿ�d���ȑ�i�j��8�^|�S+��̾���]�������̾S+�`   `   h�+��eT��6�����������?����&��'������?鿳��������6���eT�f�+��� \����������龍��!\�����`   `   ��A�f�h�9�������[ǿ�?�pW���nW��?鿰[ǿ����	9��f�h���A��@'�����;���@�������@'�`   `   8�P���s��a������������ٿگ�ݯ运�ٿ���������a����s�7�P�b|9�UM0�?�1���7�;�<�8�<���7�B�1�UM0�a|9�`   `   ۯU���s�	9�������d��|�����ſ|����d������	9����s�ݯU�{�C�$@��LI�d�X���f��Xl���f�d�X��LI�$@�{�C�`   `   8�P�i�h��6���ȑ��͝�A¤�>¤��͝��ȑ��6��f�h�7�P�{�C�@�E�z�V���p��x�����������x����p�x�V�A�E�z�C�`   `   ��A��eT�q�j������С�������i�j��eT���A�b|9�$@�z�V���y�:��JU���+��GU��:����y�z�V�$@�b|9�`   `   h�+��8�3�H�ƇV��F^��F^���V�7�H��8�f�+��@'�UM0��LI���p�:����(9��)9����9����p��LI�UM0��@'�`   `   `|����	�#�P�+�zr.�P�+�
�#����^|�����?�1�d�X��x��JU��(9������(9��IU���x��g�X�?�1�����`   `   �e�T��א��,�,�ސ��K���e�S+� \������7���f������+��)9��(9���+��������f���7���!\��K+�`   `   R���޻��쿾����쿾޻�_���ꂼ���̾���;��;�<��Xl�����GU����IU�������Xl�;�<�;����ﾚ�̾ꂼ�`   `   ��MN��ҋ�ҋ�WN����x���柾�������8�<���f��x��:��9���x����f�;�<�
���龺���柾x��`   `   "�N��qI��H��qI��N���[���v�A���]�����@����7�d�X���p���y���p�g�X���7�;�����i��A�����v���[�`   `   ���������}��C<%��?��kh�E�����������B�1��LI�x�V�z�V��LI�?�1�����ﾺ��A���lh��?�0<%�`   `   ��r׽���N��6���?���v��柾��̾!\����UM0�$@�A�E�$@�UM0���!\����̾�柾��v��?�H���N��`   `   ӝ��ĝ���ʽ�N��C<%���[�x��䂼�S+����@'�a|9�{�C�z�C�b|9��@'���K+�邼�x����[�0<%��N����ʽ`   `   �Nǽ��ؽ�w��=3�z�s�0���ؾ]�	��)���F��_�\!o�b�t�\!o��_���F��)�]�	��ؾ0����s��=3��w���ؽ`   `   ��ؽ^-���.�zs�y����R�d�З;���`�3������$��%�����4�����`�͗;�d��R�m���zs���.�^-���ؽ`   `   �w���.���s��ͫ�U���j���L�]�y�����������]�����������]�y���L��j�[���ͫ�v�s���.��w��j�`   `   �=3�zs��ͫ�0l�%%��_X��ֆ����ۢ��1�ԿAP�BP�1�Կآ������ֆ��_X�%%�6l��ͫ�zs��=3�������`   `   z�s�y���U��%%���\��H�����ӿp���Ul����Ul�r���ӿ����H����\�%%�F��y�����s���=�r,���=�`   `   0���R��j��_X��H���]��.��\��oM*���;���;�mM*�\��1���]���H���_X��j��R�0��7�w��Q��Q�?�w�`   `   �ؾd���L��ֆ����.��S�|�;��Z���f��Z�|�;�Q�.�࿎���ֆ���L�d��ؾ�:��yJ���p�uJ���:��`   `   ]�	�З;�]�y����ӿ\��|�;�`�f�cj��cj��_�f�~�;�\��ӿ���b�y�͗;�[�	��	ξK���ݏ��Ꮟ�K����	ξ`   `   �)���`�����ۢ��p���oM*��Z�cj������cj���Z�oM*�r���ۢ��������`��)�s ��c˾T�������T����c˾s �`   `   ��F�3����1�ԿUl���;���f�cj��cj����f���;�Tl�1�Կ�4�����F�����\���Ծ�Qž�Qž�Ծ�\�����`   `   �_��������AP������;��Z�_�f��Z���;����AP㿻�������_�,�0�j��ض�����E�羐��ض��g��,�0�`   `   \!o�$���]��BP�Ul�mM*�|�;�~�;�oM*�Tl�AP��]��%��Z!o���B��$����I��v	��v	�G�����$���B�`   `   b�t�%������1�Կr���\��Q�\��s���1�Կ����%��c�t��{L�Vk1�:�#���&L �� �&L ���:�#�Wk1��{L�`   `   \!o�����آ��ӿ1��.��ӿۢ������Z!o��{L��6���,�_.�=�3��Q8��Q8�@�3�].���,��6��{L�`   `   �_�4��������������]������������4����_���B�Vk1���,��13���>��I�RN��I���>��13���,�Vk1���B�`   `   ��F���`�]�y��ֆ��H���H���ֆ�b�y���`���F�,�0��$�:�#�_.���>�5+P���Z���Z�8+P���>�].�9�#��$�/�0�`   `   �)�͗;���L��_X���\��_X���L�͗;��)����j�������=�3��I���Z��a���Z��I�=�3������g�����`   `   ]�	�d��j�%%�%%��j�d�[�	�s ��\��ض��I�&L ��Q8�RN���Z���Z�PN��Q8�%L �G�޶���\��n �`   `   �ؾ�R�[��7l�F���R��ؾ�	ξ�c˾�Ծ����v	�� ��Q8��I�8+P��I��Q8�� ��v	�����Ծ�c˾�	ξ`   `   0��m����ͫ��ͫ�y���0���:��L���T����QžE���v	�&L �@�3���>���>�=�3�%L ��v	�K�羉QžJ���K����:��`   `   ��s�zs�w�s�zs���s�8�w�yJ��ݏ�������Qž���G���].��13�].���G���쾉Qž����ݏ��mJ��8�w�`   `   �=3���.���.��=3���=��Q��p�Ꮟ�T����Ծض�����:�#���,���,�9�#����޶���ԾJ���ݏ����p��Q�o�=�`   `   �w�^-��w����r,��Q�uJ��K����c˾�\��g���$�Wk1��6�Vk1��$�g���\���c˾K���mJ���Q��,����`   `   ��ؽ��ؽ�j������=�?�w��:���	ξs ����,�0���B��{L��{L���B�/�0����n ��	ξ�:��8�w�o�=�����j�`   `   �v�k(������Q�b���)�������� ���D�2ef�mՀ�ɉ��쌿ɉ�jՀ�2ef���D�� �����)���t����Q����k(��`   `   k(���P�[�M���e�Ǿ��>R2��s_��m�������`���`���������m���s_�ER2� ��W�Ǿ骏�p�M��P�S(��`   `   ���[�M�ԁ���4;���L@��v�a���i��e�Ϳ���;뿗�e�Ϳ�i��a���v��L@����4;́��[�M����U��`   `   �Q����4;_����G�<�������̿�+���o���"���"��o��+���̿���:�����G�b��
5;骏��Q� +�+�`   `   b���e�Ǿ����G�s9�����j࿥���T;���Z�3�f���Z��T;����f࿘��x9����G���e�Ǿl�����X��UC���X�`   `   )������L@�<��������?r!��Z��b��0H��/H���b���Z�Ar!��翔��:����L@� ��#���R_���Oh��Oh�V_��`   `   ����>R2��v����j�?r!���e�p���B~��>ɼ�C~��p�����e�?r!�m࿂���v�>R2�����Mc���ȍ�=���ȍ�Mc��`   `   � ��s_�a���̿����Z�p������,���+������p����Z�����̿a���s_�� �ї�$���w1��{1��#���ʗ�`   `   ��D��m���i���+���T;��b��B~��,���l���,���A~���b���T;��+���i���m����D����<�վ�έ�l)���έ�C�վ���`   `   1ef�
���e�Ϳ�o���Z�0H��>ɼ�+���,���>ɼ�/H����Z��o�h�Ϳ���.ef�'d*�����V�̾O��K��P�̾����*d*�`   `   mՀ����㿋�"�3�f�/H��C~�����A~��/H��6�f���"�����nՀ��PC�K���q���ξ��ľ��ξ�q�H���PC�`   `   ɉ�`����;뿌�"���Z��b��p���p����b����Z���"��;�`���~ɉ�V��&��8������ھ��ھ����8��&�V�`   `   �쌿`����㿚o��T;��Z���e��Z��T;��o���`����쌿M9`�"�2�l����O�����O����l��$�2�M9`�`   `   ɉ���e�Ϳ�+�����Ar!�?r!�����+��h�Ϳ��~ɉ�M9`�e�6�3���#�����U��U�����#�1��e�6�M9`�`   `   jՀ�����i���̿f���m��̿�i�����nՀ�V�"�2�3���h���	�>R	���	�8R	���	��h�3��#�2�V�`   `   2ef��m��a��������������a���m��/ef��PC��&�m���#���	��Q�f��i���Q���	��#�l���&��PC�`   `   ��D��s_��v�:���y9��:����v��s_���D�'d*�K���8������>R	�f�����f��<R	�������8�H��'d*�`   `   � �ER2��L@���G���G��L@�>R2�� ���������q��O��U���	�i��f����	��U�N�򾭞꾕q������`   `   ���� ����c���� ������ї�<�վV�̾��ξ��ھ����U�8R	��Q�<R	��U������ھ�ξV�̾H�վї�`   `   )���W�Ǿ�4;
5;e�Ǿ#���Mc��$����έ�O����ľ��ھO������	���	����N����ھ��ľK���έ�$���[c��`   `   t���ꪏ�΁��ꪏ�l���R_���ȍ�w1��l)��K����ξ������#��h��#�������ξK��{)��w1���ȍ�R_��`   `   �Q�p�M�[�M��Q���X��Oh�=��{1���έ�P�̾�q��8�m��1��3��l���8��q�V�̾�έ�w1��K���Oh���X�`   `   ����P���� +��UC��Oh��ȍ�$���C�վ����I���&�$�2�e�6�#�2��&�H������H�վ$����ȍ��Oh��UC� +�`   `   k(��S(��U��+���X�V_��Mc��ʗ澻��*d*��PC�V�N9`�M9`�V��PC�'d*����ї�[c��R_����X� +�j��`   `   �8��E�J3��m��Р��+پ���*K7�`�����'��㕜�CS��㕜�'������`�*K7�����+پѠ��m�43��E�`   `   �E�V�.���j��A��B��%��0�M�`��P���].��`Mǿj
Կj
ԿbMǿ^.��M����_��8�M�)��3���A��ƹj�T�.�tE�`   `   J3���j�����J��8�%��x^�#���j����ؿ�3����x������3���ؿ�j��!���x^�<�%�J�쾑�����j�Z3�Q� �`   `   �m��A��J��a�(���g��y���?Ŀ�o�7�(�i�N�,�e�-�e�i�N�5�(��o��?Ŀ�y���g�e�(�W���A���m���@���@�`   `   �Р�B��8�%���g�;ښ��Bп�����M�A���4;���q��4;��A�����M����Bп@ښ���g�/�%�B��
Ѡ�Bzs�u(Z�Bzs�`   `   �+پ%���x^��y���Bп(%��dd��Ş�w����c���c��v����Ş��dd�(%��Bп�y���x^�)���+پ:����P���P��>���`   `   ���0�M�#���?Ŀ����dd�ǧ����� ���
� �����ǧ��dd�����?Ŀ"��0�M������ʾ� ������� ����ʾ`   `   *K7�`���j���o���M��Ş������r
�aX�aX��r
������Ş���M��o��j���_��'K7��� ��0���
���
���0���� �`   `   `�P�����ؿ7�(�A���w��� �aX���"�aX� �w���A���7�(���ؿP���	`�v�=��J�����J��E��v�`   `   ����].���3�i�N�4;���c����
�aX�aX���
��c��3;��i�N��3�^.������ӯ=�`���cо�౾�౾�cо`��֯=�`   `   '��`Mǿ���,�e��q���c�� ��r
� ��c���q��,�e����`Mǿ'����X��O�6��þ�Z����þ6�O���X�`   `   㕜�j
Կx��,�e�4;��v�����������w���3;��,�e�y��j
Կᕜ�!�l�hv0�(���ؾ"J��J���ؾ,��hv0��l�`   `   CS��j
Կ���i�N�A����Ş�ǧ��Ş�A���i�N����j
ԿDS����w���<�����~�D�̾]yþD�̾�~������<���w�`   `   㕜�bMǿ�3�5�(���M��dd��dd���M�7�(��3�`Mǿ╜���w��@�8/�%����ؾbʾiʾ�ؾ!���6/��@���w�`   `   '��^.����ؿ�o���(%�����o���ؿ^.��'��!�l���<�8/�A����޾q�ϾU�˾c�Ͼ��޾A��8/���<�!�l�`   `   ����M����j���?Ŀ�Bп�Bп�?Ŀ�j��P���������X�hv0����%�����޾�^ҾI�;O�;�^Ҿ��޾!������hv0���X�`   `   `��_��!���y��@ښ��y��"���_��	`�ӯ=��O�(���~��ؾq�ϾI�;LO;I�;m�Ͼ�ؾ�~�(���O�ӯ=�`   `   *K7�8�M��x^��g���g��x^�0�M�'K7�v�`��6���ؾD�̾bʾU�˾O�;I�;R�˾iʾB�̾�ؾ>��`��o�`   `   ���)��<�%�e�(�/�%�)������� �=���cо��þ#J��]yþiʾc�Ͼ�^Ҿm�ϾiʾXyþ"J����þ�cоK���� �`   `   �+پ3��K��W��B�往+پ��ʾ�0��J���౾�Z��J��D�̾�ؾ��޾��޾�ؾB�̾"J���Z���౾J���0��͆ʾ`   `   Ѡ��A�������A��
Ѡ�:���� ���
������౾��þ�ؾ�~�!���A��!����~��ؾ��þ�౾-����
��� ��:���`   `   �m�ƹj���j��m�Bzs��P�������
��J���cо6��,�����6/�8/����(��>���cоJ���
�������P��#zs�`   `   43�T�.�Z3���@�v(Z��P��� ���0��E��`���O�hv0���<��@���<�hv0��O�`��K���0��� ���P���(Z���@�`   `   �E�tE�Q� ���@�Bzs�>�����ʾ�� �v�֯=���X��l���w���w�!�l���X�ӯ=�o��� �͆ʾ:���#zs���@�j� �`   `   NZ��k��SD� ������E-ﾠj�>J���v��⏿��������`�������݃���⏿��v�>J��j�E-ﾘ��� ���SD��k�`   `   �k��?� ��*!��Y���-���c�@
������˿�翃����������˿���>
���c��-�I��&!��-���?��k�`   `   �SD� ���ض�.=�j(8�D�v�E���ɿ�j{ ��9��xC��9�j{ ���ɿ�D��D�v�o(8�.=��ض� ���SD��10�`   `    ��*!��.=��;�Ye���թ��U������W��"���������"����W�����U心թ�Ue����;�5=�&!�����g�R�j�R�`   `   ����Y��j(8�Ye�����H����8��ą�7ذ�L`���y��L`��8ذ��ą��8�H������Ye��`(8�Y������΄�Pm�΄�`   `   E-��-�D�v��թ�H���#B��H������A��������A�������H��#B�C����թ�K�v��-�=-�)&��b���a���-&��`   `   �j���c�E���U��8��H������P���1+�i�4��1+�P�������H���8��U� E����c��j�;�ܾ����������;�ܾ`   `   >J�@
���ɿ����ą�����P���n4��HH��HH��n4�P�������ą�����ɿ>
��>J����6˾x{��|{���6˾���`   `   ��v�������W�7ذ�A���1+��HH�N�R��HH��1+�A��8ذ���W�������v���-��&��'��8���'���&����-�`   `   �⏿�˿j{ ��"��L`�����i�4��HH��HH�j�4����K`���"��k{ ��˿�⏿��N�&a�m�ؾ�봾�봾f�ؾ%a���N�`   `   �������9�����y������1+��n4��1+���� z������9���ს���k��
)�CW���Iþ��JþCW���
)���k�`   `   ���������xC����L`��A��P��P��A��K`������xC����������ŀ��<�2,	�ĶӾ�u���u����Ӿ5,	��<��ŀ�`   `   `��������9��"��8ذ�������������8ذ��"���9�����a���������H�7"�����ռ������ռ����7"���H�����`   `   ������j{ ���W��ą��H���H���ą���W�k{ �����������&M�)����#Sþ��� ���*Sþ���	)�&M�����`   `   ݃���˿�����8�#B��8������˿ს��ŀ���H�)�&���VǾ�^��	&���^���VǾ.��)���H��ŀ�`   `   �⏿����ɿ�U�H���C����U��ɿ����⏿��k��<�7"�����VǾVⰾ��������]ⰾ�VǾ���6"��<���k�`   `   ��v�>
���D���թ�����թ� E��>
����v���N��
)�2,	����#Sþ�^�������֣������^��#Sþ���2,	��
)���N�`   `   >J��c�D�v�Ue��Ye��K�v���c�>J���-�&a�CW��ĶӾ�ռ����	&����������&�� ����ռ���ӾKW��%a���-�`   `   �j��-�o(8���;�`(8��-��j����&��n�ؾ�Iþ�u������ ����^��]ⰾ�^�� ���񺰾�u���Iþn�ؾ�&����`   `   E-�I��/=�5=�Z��>-�<�ܾ�6˾'���봾���u���ռ�*Sþ�VǾ�VǾ#Sþ�ռ��u�����봾'���6˾L�ܾ`   `   ����&!���ض�&!������*&�����x{��8����봾Jþ��Ӿ������.���������Ӿ�Iþ�봾J���x{�����*&��`   `    ��-�� �����΄�b�������|{��'��g�ؾCW��6,	�7"�
)�)�6"�2,	�KW��n�ؾ'��x{������a����̈́�`   `   �SD��?��SD�h�R�Pm�a�������6˾�&��&a��
)��<���H�&M���H��<��
)�&a��&���6˾���a���8Pm�h�R�`   `   �k��k��10�j�R�΄�.&��<�ܾ�����-���N���k��ŀ����������ŀ���k���N���-���L�ܾ)&���̈́�h�R�20�`   `   t���(���O�x���v�����Q(��V�t���aܘ�T���1ں��2��1ں�Q���aܘ�y����V�Q(�������w�����O��(�`   `   �(�N�J�]���>4��4 ���8���q�T<��踿�p޿��
7�
7����p޿	踿R<����q���8�+ �:4��k���K�J��(�`   `   ��O�]���`#¾~��)D���'����ݿ��[�8�&�W�Wc�%�W�[�8�����ݿ$�����.D�~��V#¾]�����O��':�`   `   w���>4��~��G�G��������b���>8���|�J����`���`��J�����|�>8�g�������K�G����94��o����^��^�`   `   v��4 �)D������&���
�ӍV�[_��{e���r��YA��r��|e��[_��ЍV��
��&������D�4 ����$���	z�$��`   `   �����8�������
��.b����-���X���*���*��X��-�����.b��
��������8����I���K��J��M���`   `   Q(���q�'���b���ӍV���m�ʧ*�\�G��dR�]�G�ʧ*�l���ԍV�b���%�����q�Q(�:��jZ���Ŝ�hZ��:��`   `   �V�S<���ݿ>8�[_���-��ʧ*�#UR��i��i�#UR�˧*��-��Y_��>8��ݿR<���V����.վVy��[y���.վ��`   `   t���踿����|�{e���X�\�G��i��tu��i�\�G��X�|e����|���踿w�����7����Bľ�����Bľ����7�`   `   `ܘ��p޿[�8�J����r����*��dR��i��i��dR���*��r��J���\�8��p޿^ܘ���Z��x�`�߾��������Y�߾�x���Z�`   `   T�����&�W��`��YA���*�]�G�#UR�\�G���*�ZA��`��$�W���U���	y�1�t���s�žR峾~�žt���1�	y�`   `   1ں�
7�Wc��`���r���X�ʧ*�˧*��X��r���`��Wc�
7�/ں�އ���D���P�Ծ�"���"��K�Ծ����D�އ�`   `   �2��
7�%�W�J���|e���-��l��-��|e��J���$�W�
7��2��_���a�Q�$�Q�⾴���&驾����O��$�c�Q�_���`   `   1ں���[�8���|�[_������Y_����|�\�8���/ں�_���i�V��3�"���𻾙����������3�h�V�^���`   `   Q����p޿���>8�ЍV��.b�ԍV�>8����p޿U���އ�a�Q��3��M�%���L��Ȋ���K��%���N��3�c�Q�އ�`   `   aܘ�	踿�ݿg����
��
�b����ݿ踿_ܘ�
y���D�$�"��%���\좾��c좾"�����$���D�y�`   `   y���R<��$�������&�����%���R<��x�����Z�1���Q����L��������L����X�⾂�1���Z�`   `   �V���q������������q��V���7��x�t���P�Ծ�������Ȋ����Ŋ���������L�Ծ}����x���7�`   `   Q(���8�.D�K�G�D���8�Q(�����`�߾s�ž�"��&驾����K��c좾L�����!驾�"��n�ž`�߾����`   `   ���+ �~�����4 ����:�龅.վ�Bľ����R峾�"��������&���"����𻾲����"��[峾�����Bľ�.վL��`   `   ���:4��V#¾:4�����I���jZ��Wy����������~�žL�ԾO����N���X��L�Ծn�ž�������Wy��ZZ��I���`   `   x���k���]���o���$��K���Ŝ�[y���BľY�߾t�����$��3��3�$���}���`�߾�BľWy���Ŝ�J��$��`   `   ��O�K�J���O��^��	z�J��hZ���.վ���x�1���D�d�Q�h�V�c�Q���D�1��x����.վZZ��J��
z��^�`   `   �(��(��':��^�$��N���:������7���Z�
y�އ�_���^���އ�y���Z���7���L��I���$���^��':�`   `   '��N�+��qS�Z!�������z���+�q	[��U��������𪿿eUſ謹��������U��q	[���+��z�����Z!���qS�N�+�`   `   N�+���N��M��mľ��	���<��v�ʄ��ͽ�v�応�U�U���w��ͽ�Ȅ���v���<���	�iľ�M����N�=�+�`   `   �qS��M���ƾV��k9H��΅��ŭ�������A���b�[bo���b���A�������ŭ��΅�p9H�V���ƾ�M���qS���=�`   `   Z!��mľV��I4L�z��	�����mIA��,���k��Q7��Q7���k���,��nIA����	���y��M4L�]��iľR!����b���b�`   `   ������	�j9H�z���g��u��A�a�>4�����
�Jj	��
���>4��>�a�u���g��z��`9H���	�����������~�����`   `   �z���<��΅�	��u��s^n��ݹ����v�!���3���3�v�!�����ݹ�s^n�s��	���΅���<��z�c����������g��`   `   ��+��v��ŭ����A�a��ݹ��F	���3��*R��<]��*R���3��F	��ݹ�C�a�����ŭ��v���+�M���R���G���R��M��`   `   q	[�ʄ�����mIA�>4�������3��1]�@u�@u��1]���3����=4��nIA����Ȅ��m	[�ڔ���ؾg��k����ؾה�`   `   �U��ͽ�~��,����v�!��*R�@u�t��@u��*R�v�!����,��|�ͽ��U���|;�$B���ƾ&�����ƾ(B��|;�`   `   ���v����A��k���
���3��<]�@u�@u��<]���3��
��k����A�w�忻��|�^�'���⾰����������&���^�`   `   �������b�Q7��Jj	���3��*R��1]��*R���3�Kj	�Q7����b�������}��4�� ��Ǿ襴��Ǿ� ��4��}�`   `   謹�U�[bo�Q7���
�v�!���3���3�v�!��
�Q7��]bo�U���vf���H����]�վG�@�Y�վ����H�uf��`   `   eUſU���b��k��������F	�������k����b�U�gUſ����ZYU�����\����<[������\㾆��]YU�����`   `   謹�����A��,��>4���ݹ��ݹ�=4���,����A�����������Y�U����L��Q_��Y_��L����S����Y�����`   `   ���w�忀�nIA�>�a�s^n�C�a�nIA�|�w�����vf��ZYU�U����ü����:�������ü���U��\YU�vf��`   `   ���ͽ���俳��u��s��������ͽ�����}��H������ü�P=��x^��^��W=���ü������H��}�`   `   �U��Ȅ���ŭ�	���g��	���ŭ�Ȅ���U��|�^��4�����\�L�����x^��hȌ�x^�����L���\㾢���4�|�^�`   `   q	[��v��΅��y��z���΅��v�m	[��|;�'�� �]�վ���R_��:���^��x^��7���Y_�����Y�վ� �&��|;�`   `   ��+���<�p9H�M4L�`9H���<���+�ڔ�$B���⾶ǾG�<[��Y_�����W=�����Y_��7[��G󳾱Ǿ���,B�ڔ�`   `   �z���	�V��]����	��z�M���ؾ��ƾ����襴�@����L���ü��ü�L�����G�񥴾������ƾ��ؾ_��`   `   ����iľ�ƾiľ����c���R��g��&��������ǾY�վ�\��������\�Y�վ�Ǿ����9���g���R��c��`   `   Z!���M���M��R!�����������G��k����ƾ���� �������S��U��������� ������ƾg��
H������괎�`   `   �qS���N��qS���b���~������R����ؾ(B�&��4��H�]YU���Y�\YU��H��4�&�,B���ؾ�R�������~���b�`   `   N�+�=�+���=���b�����g��M��ה��|;���^��}�uf����������vf���}�|�^��|;�ڔ�_��c��괎���b�Ř=�`   `   t���(���O�w���v�����Q(��V�t���aܘ�T���1ں��2��1ں�Q���aܘ�y����V�Q(�������w�����O��(�`   `   �(�N�J�]���>4��4 ���8���q�T<��踿�p޿��
7�
7����p޿	踿R<����q���8�+ �:4��k���K�J��(�`   `   ��O�]���`#¾~��)D���'����ݿ��[�8�&�W�Wc�%�W�[�8�����ݿ$�����.D�~��V#¾]�����O��':�`   `   w���>4��~��G�G��������b���>8���|�J����`���`��J�����|�>8�g�������K�G����94��o����^��^�`   `   v��4 �)D������&���
�ӍV�[_��{e���r��YA��r��|e��[_��ЍV��
��&������D�4 ����$���	z�$��`   `   �����8�������
��.b����-���X���*���*��X��-�����.b��
��������8����I���K��J��M���`   `   Q(���q�'���b���ӍV���m�ʧ*�\�G��dR�]�G�ʧ*�l���ԍV�b���%�����q�Q(�:��jZ���Ŝ�hZ��:��`   `   �V�S<���ݿ>8�[_���-��ʧ*�#UR��i��i�#UR�˧*��-��Y_��>8��ݿR<���V����.վVy��[y���.վ��`   `   t���踿����|�{e���X�\�G��i��tu��i�\�G��X�|e����|���踿w�����7����Bľ�����Bľ����7�`   `   `ܘ��p޿[�8�J����r����*��dR��i��i��dR���*��r��J���\�8��p޿^ܘ���Z��x�`�߾��������Y�߾�x���Z�`   `   T�����&�W��`��YA���*�]�G�#UR�\�G���*�ZA��`��$�W���U���	y�1�t���s�žR峾~�žt���1�	y�`   `   1ں�
7�Wc��`���r���X�ʧ*�˧*��X��r���`��Wc�
7�/ں�އ���D���P�Ծ�"���"��L�Ծ����D�އ�`   `   �2��
7�%�W�J���|e���-��l��-��|e��J���$�W�
7��2��_���a�Q�$�Q�⾴���&驾����O��$�c�Q�_���`   `   1ں���[�8���|�[_������Y_����|�\�8���/ں�_���i�V��3�"���𻾙����������3�h�V�^���`   `   Q����p޿���>8�ЍV��.b�ԍV�>8����p޿U���އ�a�Q��3��M�%���L��Ȋ���K��%���N��3�c�Q�އ�`   `   aܘ�	踿�ݿg����
��
�b����ݿ踿_ܘ�
y���D�$�"��%���\좾��c좾"�����$���D�y�`   `   y���R<��$�������&�����%���R<��x�����Z�1���Q����L��������L����X�⾂�1���Z�`   `   �V���q������������q��V���7��x�t���P�Ծ�������Ȋ����Ŋ���������L�Ծ}����x���7�`   `   Q(���8�.D�K�G�D���8�Q(�����`�߾s�ž�"��&驾����K��c좾L�����!驾�"��n�ž`�߾����`   `   ���+ �~�����4 ����:�龅.վ�Bľ����R峾�"��������&���"����𻾲����"��[峾�����Bľ�.վL��`   `   ���:4��V#¾:4�����I���jZ��Wy����������~�žL�ԾO����N���X��L�Ծn�ž�������Wy��ZZ��I���`   `   x���k���]���o���$��K���Ŝ�[y���BľY�߾t�����$��3��3�$���}���`�߾�BľWy���Ŝ�J��$��`   `   ��O�K�J���O��^��	z�J��hZ���.վ���x�1���D�d�Q�h�V�c�Q���D�1��x����.վZZ��J��
z��^�`   `   �(��(��':��^�$��N���:������7���Z�
y�އ�_���^���އ�y���Z���7���L��I���$���^��':�`   `   NZ��k��SD� ������E-ﾠj�>J���v��⏿��������`�������݃���⏿��v�>J��j�E-ﾘ��� ���SD��k�`   `   �k��?� ��*!��Y���-���c�@
������˿�翃����������˿���>
���c��-�I��&!��-���?��k�`   `   �SD����ض�.=�j(8�D�v�E���ɿ�j{ ��9��xC��9�j{ ���ɿ�D��D�v�o(8�.=��ض� ���SD��10�`   `    ��*!��.=��;�Ye���թ��U������W��"���������"����W�����U心թ�Ue����;�5=�&!�����g�R�j�R�`   `   ����Y��j(8�Ye�����H����8��ą�7ذ�L`���y��L`��8ذ��ą��8�H������Ye��`(8�Y������΄�Pm�΄�`   `   E-��-�D�v��թ�H���#B��H������A��������A�������H��#B�C����թ�K�v��-�=-�)&��b���a���-&��`   `   �j���c�E���U��8��H������P���1+�i�4��1+�P�������H���8��U� E����c��j�;�ܾ����������;�ܾ`   `   >J�@
���ɿ����ą�����P���n4��HH��HH��n4�P�������ą�����ɿ>
��>J����6˾x{��|{���6˾���`   `   ��v�������W�7ذ�A���1+��HH�N�R��HH��1+�A��8ذ���W�������v���-��&��'��8���'���&����-�`   `   �⏿�˿j{ ��"��L`�����i�4��HH��HH�j�4����K`���"��k{ ��˿�⏿��N�&a�m�ؾ�봾�봾f�ؾ%a���N�`   `   �������9�����y������1+��n4��1+���� z������9���ს���k��
)�CW���Iþ��JþCW���
)���k�`   `   ���������xC����L`��A��P��P��A��K`������xC����������ŀ��<�2,	�ĶӾ�u���u����Ӿ5,	��<��ŀ�`   `   `��������9��"��8ذ�������������8ذ��"���9�����a���������H�7"�����ռ������ռ����7"���H�����`   `   ������j{ ���W��ą��H���H���ą���W�k{ �����������&M�)����#Sþ��� ���*Sþ���	)�&M�����`   `   ݃���˿�����8�#B��8������˿ს��ŀ���H�)�&���VǾ�^��	&���^���VǾ.��)���H��ŀ�`   `   �⏿����ɿ�U�H���C����U��ɿ����⏿��k��<�7"�����VǾVⰾ��������]ⰾ�VǾ���6"��<���k�`   `   ��v�>
���D���թ�����թ� E��>
����v���N��
)�2,	����#Sþ�^�������֣������^��#Sþ���2,	��
)���N�`   `   >J��c�D�v�Ue��Ye��K�v���c�>J���-�&a�CW��ĶӾ�ռ����	&����������&�� ����ռ���ӾKW��&a���-�`   `   �j��-�o(8���;�`(8��-��j����&��n�ؾ�Iþ�u������ ����^��]ⰾ�^�� ���񺰾�u���Iþn�ؾ�&����`   `   E-�I��/=�5=�Z��>-�<�ܾ�6˾'���봾���u���ռ�*Sþ�VǾ�VǾ#Sþ�ռ��u�����봾'���6˾L�ܾ`   `   ����&!���ض�&!������*&�����x{��8����봾Jþ��Ӿ������.���������Ӿ�Iþ�봾J���x{�����*&��`   `    ��-�� �����΄�b�������|{��'��g�ؾCW��6,	�7"�
)�)�6"�2,	�KW��n�ؾ'��x{������a����̈́�`   `   �SD��?��SD�h�R�Pm�a�������6˾�&��&a��
)��<���H�&M���H��<��
)�&a��&���6˾���a���8Pm�h�R�`   `   �k��k��10�j�R�΄�.&��<�ܾ�����-���N���k��ŀ����������ŀ���k���N���-���L�ܾ)&���̈́�h�R�20�`   `   �8��E�J3��m��Р��+پ���*K7�`�����'��㕜�CS��㕜�'������`�*K7�����+پѠ��m�43��E�`   `   �E�V�.���j��A��B��%��0�M�`��P���].��`Mǿj
Կj
ԿbMǿ^.��M����_��8�M�)��3���A��Źj�T�.�tE�`   `   J3���j�����J��8�%��x^�#���j����ؿ�3����x������3���ؿ�j��!���x^�<�%�J�쾑�����j�Z3�Q� �`   `   �m��A��J��a�(���g��y���?Ŀ�o�7�(�i�N�,�e�-�e�i�N�5�(��o��?Ŀ�y���g�e�(�W���A���m���@���@�`   `   �Р�B��8�%���g�;ښ��Bп�����M�A���4;���q��4;��A�����M����Bп@ښ���g�/�%�B��
Ѡ�Bzs�u(Z�Bzs�`   `   �+پ%���x^��y���Bп(%��dd��Ş�w����c���c��v����Ş��dd�(%��Bп�y���x^�)���+پ:����P���P��>���`   `   ���0�M�#���?Ŀ����dd�ǧ����� ���
� �����ǧ��dd�����?Ŀ"��0�M������ʾ� ������� ����ʾ`   `   *K7�`���j���o���M��Ş������r
�aX�aX��r
������Ş���M��o��j���_��'K7��� ��0���
���
���0���� �`   `   `�P�����ؿ7�(�A���w��� �aX���"�aX� �w���A���7�(���ؿP���	`�v�=��J�����J��E��v�`   `   ����].���3�i�N�4;���c����
�aX�aX���
��c��3;��i�N��3�^.������ӯ=�`���cо�౾�౾�cо`��֯=�`   `   '��`Mǿ���,�e��q���c�� ��r
� ��c���q��,�e����`Mǿ'����X��O�6��þ�Z����þ6�O���X�`   `   㕜�j
Կx��-�e�4;��v�����������w���3;��,�e�y��j
Կᕜ�!�l�hv0�(���ؾ"J��J���ؾ,��hv0��l�`   `   CS��j
Կ���i�N�A����Ş�ǧ��Ş�A���i�N����j
ԿDS����w���<�����~�D�̾]yþD�̾�~������<���w�`   `   㕜�bMǿ�3�5�(���M��dd��dd���M�7�(��3�`Mǿ╜���w��@�8/�%����ؾbʾiʾ�ؾ!���6/��@���w�`   `   '��^.����ؿ�o���(%�����o���ؿ^.��'��!�l���<�8/�A����޾q�ϾU�˾c�Ͼ��޾A��8/���<�!�l�`   `   ����M����j���?Ŀ�Bп�Bп�?Ŀ�j��P���������X�hv0����%�����޾�^ҾI�;O�;�^Ҿ��޾!������hv0���X�`   `   `��_��!���y��@ښ��y��"���_��	`�ӯ=��O�(���~��ؾq�ϾI�;MO;I�;m�Ͼ�ؾ�~�(���O�ӯ=�`   `   *K7�8�M��x^��g���g��x^�0�M�'K7�v�`��6���ؾD�̾bʾU�˾O�;I�;R�˾iʾB�̾�ؾ>��`��o�`   `   ���)��<�%�e�(�/�%�)������� �=���cо��þ#J��]yþiʾc�Ͼ�^Ҿm�ϾiʾXyþ"J����þ�cоK���� �`   `   �+پ3��K��W��B�往+پ��ʾ�0��J���౾�Z��J��D�̾�ؾ��޾��޾�ؾB�̾#J���Z���౾J���0��͆ʾ`   `   Ѡ��A�������A��
Ѡ�:���� ���
������౾��þ�ؾ�~�!���A��!����~��ؾ��þ�౾-����
��� ��:���`   `   �m�ƹj���j��m�Bzs��P�������
��J���cо6��,�����6/�8/����(��>���cоJ���
�������P��#zs�`   `   43�T�.�Z3���@�v(Z��P��� ���0��E��`���O�hv0���<��@���<�hv0��O�`��K���0��� ���P���(Z���@�`   `   �E�tE�Q� ���@�Bzs�>�����ʾ�� �v�֯=���X��l���w���w�!�l���X�ӯ=�o��� �͆ʾ:���#zs���@�j� �`   `   �v�k(������Q�b���)�������� ���D�2ef�mՀ�ɉ��쌿ɉ�jՀ�2ef���D�� �����)���t����Q����k(��`   `   k(���P�[�M���e�Ǿ��>R2��s_��m�������`���`���������m���s_�ER2� ��W�Ǿ骏�p�M��P�S(��`   `   ���[�M�ԁ���4;���L@��v�a���i��e�Ϳ���;뿗�e�Ϳ�i��a���v��L@����4;́��[�M����U��`   `   �Q����4;_����G�<�������̿�+���o���"���"��o��+���̿���:�����G�b��
5;骏��Q� +�+�`   `   b���e�Ǿ����G�s9�����j࿥���T;���Z�3�f���Z��T;����f࿘��x9����G���e�Ǿl�����X��UC���X�`   `   )������L@�<��������?r!��Z��b��0H��/H���b���Z�Ar!��翔��:����L@� ��#���R_���Oh��Oh�V_��`   `   ����>R2��v����j�?r!���e�p���B~��>ɼ�C~��p�����e�?r!�m࿂���v�>R2�����Mc���ȍ�=���ȍ�Mc��`   `   � ��s_�a���̿����Z�p������,���+������p����Z�����̿a���s_�� �ї�$���w1��{1��#���ʗ�`   `   ��D��m���i���+���T;��b��B~��,���l���,���A~���b���T;��+���i���m����D����<�վ�έ�l)���έ�C�վ���`   `   1ef�
���e�Ϳ�o���Z�0H��>ɼ�+���,���>ɼ�/H����Z��o�h�Ϳ���.ef�'d*�����V�̾O��K��P�̾����*d*�`   `   mՀ����㿋�"�3�f�/H��C~�����A~��/H��6�f���"�����nՀ��PC�K���q���ξ��ľ��ξ�q�H���PC�`   `   ɉ�`����;뿌�"���Z��b��p���p����b����Z���"��;�`���~ɉ�V��&��8������ھ��ھ����8��&�V�`   `   �쌿`����㿚o��T;��Z���e��Z��T;��o���`����쌿M9`�"�2�l����O�����O����l��$�2�M9`�`   `   ɉ���e�Ϳ�+�����Ar!�?r!�����+��h�Ϳ��~ɉ�M9`�e�6�3���#�����U��U�����#�1��e�6�M9`�`   `   jՀ�����i���̿f���m��̿�i�����nՀ�V�"�2�3���h���	�>R	���	�8R	���	��h�3��#�2�V�`   `   2ef��m��a��������������a���m��/ef��PC��&�m���#���	��Q�f��i���Q���	��#�l���&��PC�`   `   ��D��s_��v�:���y9��:����v��s_���D�'d*�K���8������>R	�f�����f��<R	�������8�H��'d*�`   `   � �ER2��L@���G���G��L@�>R2�� ���������q��O��U���	�j��f����	��U�N�򾭞꾕q������`   `   ���� ����c���� ������ї�<�վV�̾��ξ��ھ����U�8R	��Q�<R	��U������ھ�ξV�̾H�վї�`   `   )���W�Ǿ�4;
5;e�Ǿ#���Mc��$����έ�O����ľ��ھO������	���	����N����ھ��ľK���έ�$���[c��`   `   t���ꪏ�΁��ꪏ�l���R_���ȍ�w1��l)��K����ξ������#��h��#�������ξK��{)��w1���ȍ�R_��`   `   �Q�p�M�[�M��Q���X��Oh�=��{1���έ�P�̾�q��8�m��1��3��l���8��q�V�̾�έ�w1��K���Oh���X�`   `   ����P���� +��UC��Oh��ȍ�$���C�վ����I���&�$�2�e�6�#�2��&�H������H�վ$����ȍ��Oh��UC� +�`   `   k(��S(��U��+���X�V_��Mc��ʗ澻��*d*��PC�V�N9`�M9`�V��PC�'d*����ї�[c��R_����X� +�j��`   `   �Nǽ��ؽ�w��=3�z�s�0���ؾ]�	��)���F��_�\!o�b�t�\!o��_���F��)�]�	��ؾ0����s��=3��w���ؽ`   `   ��ؽ^-���.�zs�y����R�d�З;���`�3������$��%�����4�����`�͗;�d��R�m���zs���.�^-���ؽ`   `   �w���.���s��ͫ�U���j���L�]�y�����������]�����������]�y���L��j�[���ͫ�v�s���.��w��j�`   `   �=3�zs��ͫ�0l�%%��_X��ֆ����ۢ��1�ԿAP�BP�1�Կآ������ֆ��_X�%%�6l��ͫ�zs��=3�������`   `   z�s�y���U��%%���\��H�����ӿp���Ul����Ul�r���ӿ����H����\�%%�F��y�����s���=�r,���=�`   `   0���R��j��_X��H���]��.��\��oM*���;���;�mM*�\��1���]���H���_X��j��R�0��7�w��Q��Q�?�w�`   `   �ؾd���L��ֆ����.��S�|�;��Z���f��Z�|�;�Q�.�࿎���ֆ���L�d��ؾ�:��yJ���p�uJ���:��`   `   ]�	�З;�]�y����ӿ\��|�;�`�f�cj��cj��_�f�~�;�\��ӿ���b�y�͗;�[�	��	ξK���ݏ��Ꮟ�K����	ξ`   `   �)���`�����ۢ��p���oM*��Z�cj������cj���Z�oM*�r���ۢ��������`��)�s ��c˾T�������T����c˾s �`   `   ��F�3����1�ԿUl���;���f�cj��cj����f���;�Tl�1�Կ�4�����F�����\���Ծ�Qž�Qž�Ծ�\�����`   `   �_��������AP������;��Z�_�f��Z���;����AP㿻�������_�,�0�j��ض�����E�羐��ض��g��,�0�`   `   \!o�$���]��BP�Ul�mM*�|�;�~�;�oM*�Tl�AP��]��%��Z!o���B��$����I��v	��v	�G�����$���B�`   `   b�t�%������1�Կr���\��Q�\��s���1�Կ����%��c�t��{L�Vk1�:�#���&L �� �&L ���:�#�Wk1��{L�`   `   \!o�����آ��ӿ1��.��ӿۢ������Z!o��{L��6���,�_.�=�3��Q8��Q8�@�3�].���,��6��{L�`   `   �_�4��������������]������������4����_���B�Vk1���,��13���>��I�RN��I���>��13���,�Vk1���B�`   `   ��F���`�]�y��ֆ��H���H���ֆ�b�y���`���F�,�0��$�:�#�_.���>�5+P���Z���Z�8+P���>�].�9�#��$�/�0�`   `   �)�͗;���L��_X���\��_X���L�͗;��)����j�������=�3��I���Z��a���Z��I�=�3������g�����`   `   ]�	�d��j�%%�%%��j�d�[�	�s ��\��ض��I�&L ��Q8�RN���Z���Z�PN��Q8�%L �G�޶���\��n �`   `   �ؾ�R�[��7l�F���R��ؾ�	ξ�c˾�Ծ����v	�� ��Q8��I�8+P��I��Q8�	� ��v	�����Ծ�c˾�	ξ`   `   0��m����ͫ��ͫ�y���0���:��L���T����QžE���v	�&L �@�3���>���>�=�3�%L ��v	�K�羉QžJ���K����:��`   `   ��s�zs�w�s�zs���s�8�w�yJ��ݏ�������Qž���G���].��13�].���G���쾉Qž����ݏ��mJ��8�w�`   `   �=3���.���.��=3���=��Q��p�Ꮟ�T����Ծض�����:�#���,���,�9�#����޶���ԾJ���ݏ����p��Q�o�=�`   `   �w�^-��w����r,��Q�uJ��K����c˾�\��g���$�Wk1��6�Vk1��$�g���\���c˾K���mJ���Q��,����`   `   ��ؽ��ؽ�j������=�?�w��:���	ξs ����,�0���B��{L��{L���B�/�0����n ��	ξ�:��7�w�o�=�����j�`   `   T���ҝ���ང���N���a����e�Y|�h�+���A�8�P�ۯU�8�P���A�h�+�`|��e�R�����"�N������ҝ��`   `   ҝ��q׽����qI�WN��޻�J������8��eT�f�h���s���s�i�h��eT��8����T��޻�MN���qI����r׽ĝ��`   `   �འ���H�ҋ��쿾א���#�3�H�n�j��6��9���a��
9���6��q�j�3�H�	�#�א���쿾ҋ��H�������ʽ`   `   ����qI�ҋ����,�R�+���V����ȑ������������������ȑ���ƇV�P�+�,����ҋ��qI�|���N���N��`   `   �N�WN���쿾,�sr.��F^�����͝��d�������[ǿ�����d���͝�����F^�zr.�,��쿾WN���N�C<%�6��C<%�`   `   ��޻�֐��R�+��F^�ϡ��>¤�|�����ٿ�?��?鿎�ٿ|���A¤�С���F^�P�+�ސ��޻�
����[��?��?���[�`   `   a���J���#���V����>¤���ſگ�nW����pW�گ迼�ſ>¤������V�
�#�J��_���x����v��kh���v�x��`   `   �e쾼��3�H����͝�|���گ���'��&����ݯ�|����͝���7�H�����e�邼��柾A���E����柾䂼�`   `   Y|��8�n�j��ȑ��d����ٿnW�'��J��'��nW���ٿ�d���ȑ�i�j��8�^|�S+��̾���]�������̾S+�`   `   h�+��eT��6�����������?����&��'������?鿳��������6���eT�f�+��� \����������龍��!\�����`   `   ��A�f�h�9�������[ǿ�?�pW���nW��?鿰[ǿ����	9��f�h���A��@'�����;���@�������@'�`   `   8�P���s��a������������ٿگ�ݯ运�ٿ���������a����s�7�P�b|9�UM0�?�1���7�;�<�8�<���7�B�1�UM0�a|9�`   `   ۯU���s�	9�������d��|�����ſ|����d������	9����s�ݯU�{�C�$@��LI�d�X���f��Xl���f�d�X��LI�$@�{�C�`   `   8�P�i�h��6���ȑ��͝�A¤�>¤��͝��ȑ��6��f�h�7�P�{�C�@�E�z�V���p��x�����������x����p�x�V�A�E�z�C�`   `   ��A��eT�q�j������С�������i�j��eT���A�b|9�$@�z�V���y�:��JU���+��GU��:����y�z�V�$@�b|9�`   `   h�+��8�3�H�ƇV��F^��F^���V�7�H��8�f�+��@'�UM0��LI���p�:����(9��)9����9����p��LI�UM0��@'�`   `   `|����	�#�P�+�zr.�P�+�
�#����^|�����?�1�d�X��x��JU��(9������(9��IU���x��g�X�?�1�����`   `   �e�T��א��,�,�ސ��J���e�S+� \������7���f������+��)9��(9���+��������f���7���!\��K+�`   `   R���޻��쿾����쿾޻�_���ꂼ���̾���;��;�<��Xl�����GU����IU�������Xl�;�<�;����ﾚ�̾ꂼ�`   `   ��MN��ҋ�ҋ�WN����x���柾�������8�<���f��x��:��:���x����f�;�<�
���龺���柾x��`   `   "�N��qI��H��qI��N���[���v�A���]�����@����7�d�X���p���y���p�g�X���7�;�����i��A�����v���[�`   `   ���������}��C<%��?��kh�E�����������B�1��LI�x�V�z�V��LI�?�1�����ﾺ��A���lh��?�0<%�`   `   ��r׽���N��6���?���v��柾��̾!\����UM0�$@�A�E�$@�UM0���!\����̾�柾��v��?�H���N��`   `   ҝ��ĝ���ʽ�N��C<%���[�x��䂼�S+����@'�a|9�{�C�z�C�b|9��@'���K+�邼�x����[�0<%��N����ʽ`   `   xǃ��ܐ��˸��\��Z0�nr�����ߔо���;�P/��=�(�B��=�P/�;����ߔо����nr�0Z0��\���˸��ܐ�`   `   �ܐ�8䮽�����$�cEd�������Ⱦ�(��<���=/�Z�@���J���J�\�@��=/�9���(���Ⱦ����UEd���$���:䮽�ܐ�`   `   �˸�����o!��|_����G ɾ. ���yW8�۫N�(J]�t_b�&J]�۫N�{W8���. �G ɾ����|_��o!�����˸�;�`   `   �\����$��|_��旾1�ʾW�9�#���C���_��6t����6t���_���C�<�#�W�*�ʾ�旾�|_���$��\���ؽ�ؽ`   `   Z0�cEd����1�ʾU���i(��
M��zn�u���R���`���R���v����zn��
M��i(�[��1�ʾ���cEd�&Z0��V�6���V�`   `   nr�����G ɾW��i(��gP�S�v��&��y���x(��w(��w����&��W�v��gP��i(�W�M ɾ����ir���H��>5��>5���H�`   `   ������Ⱦ. �8�#��
M�S�v��ڎ������r��կ��r�������ڎ�S�v��
M�9�#�. ���Ⱦ����&����u��'m��u�&���`   `   ߔо�(������C��zn��&������ͥ��I��G��̥�������&���zn���C���(��ܔоVU���o��� ��� ���o��RU��`   `   ���<��yW8���_�u���y����r��I���6��I���r��y���v�����_�uW8�<�����G�{{ݾj�پR�ؾj�پ{ݾG�`   `   ;��=/�۫N��6t�R���x(��կ�G��I��կ�w(��Q����6t�ޫN��=/��:�EN�������X��X������FN�`   `   P/�Z�@�(J]��`���w(���r��̥���r��w(��c����%J]�Z�@�P/��*�a�0�na<�D9G� �K�H9G�na<�_�0��*�`   `   �=���J�t_b��R���w�����������y���Q����w_b���J��=��u?� [O��h����]b��\b�����h� [O��u?�`   `   (�B���J�&J]��6t�v����&���ڎ��&��v����6t�%J]���J�)�B��K��'e�z��P������:д����P���z���'e��K�`   `   �=�\�@�۫N���_��zn�W�v�S�v��zn���_�ޫN�Z�@��=��K��m�d%��{c����Ͽ���⿝�Ͽzc��d%���m��K�`   `   P/��=/�{W8���C��
M��gP��
M���C�uW8��=/�P/��u?��'e�d%���'��"�㿤���	����"���'��d%���'e��u?�`   `   ;�9����<�#��i(��i(�9�#���<���:��*� [O�z��{c��"�㿩J	��������J	�!��zc��z�� [O��*�`   `   ����(��. �W�[��W�. ��(�����EN�a�0��h�P�����Ͽ������' ���������ϿQ����h�_�0�EN�`   `   ߔо�ȾH ɾ*�ʾ1�ʾM ɾ��ȾݔоG����na<����������	��������	���������pa<����G�`   `   ������������旾�����������WU��{{ݾ��D9G�]b��:д��⿣���J	������9д�]b��D9G����{ݾWU��`   `   nr�UEd��|_��|_�dEd�ir�&����o��j�پ�X� �K�\b�������Ͽ"��!�㿜�Ͽ���]b��"�K��X�d�پ�o��.���`   `   0Z0���$��o!���$�&Z0���H��u�� ��R�ؾ�X�H9G����P���zc���'��zc��Q������D9G��X�[�ؾ� ���u���H�`   `   �\��������\���V��>5��'m�� ��j�پ��na<�h�z��d%��d%��z���h�pa<���d�پ� ���'m��>5��V�`   `   �˸�;䮽�˸��ؽ6���>5��u��o��{ݾ���_�0� [O��'e��m��'e� [O�_�0�����{ݾ�o���u��>5�C���ؽ`   `   �ܐ��ܐ�;��ؽ�V���H�&���RU��G�GN��*��u?��K��K��u?��*�EN�G�WU��.�����H��V��ؽP�`   `   �S��&k������Vؽ�;��MX�'P��_����������7*� �9�U?� �9��7*�������_���P���MX��;��Vؽ�����&k�`   `   �&k��Z��D���Ɇ�#�<�YO���g����ԾA�����%��\.��\.���%�	��?���Ծ�g��]O���<�Ć�R����Z���&k�`   `   ����D���n���1��Mp���E�Ⱦԓ��m,���!�+�-��2�)�-���!�o,�ԓ��C�Ⱦ���Mp��1�l��D��������ƌ�`   `   �VؽɆ��1��k�4���V�ž����b��4�&�#�6�s�>�u�>�$�6�2�&�b������S�ž/����k��1�Ć��Vؽj���g���`   `   �;�#�<��Mp�4���vrž�����S���-� �A���N��gS���N�"�A���-��S�����~rž4����Mp�#�<��;��k�� ��k�`   `   �MX�YO����V�ž�������rj2�w�J�_�\���e���e�]�\�x�J�tj2��������S�ž��]O���MX��@��4��4��@�`   `   'P���g��E�Ⱦ�����S�rj2�U�M��6d��r�d�w�"�r��6d�R�M�rj2��S�����E�Ⱦ�g��%P��?��{��ǹ�x��?��`   `   _�����Ծԓ��b����-�w�J��6d��Hw�� ��Hw��6d�x�J���-�b��ד����Ծ^����x��1ȷ��K���K��2ȷ��x��`   `   ���A�m,�4�&� �A�_�\��r���[����r�_�\�"�A�4�&�k,�A�����������B!���������`   `   �������!�#�6���N���e�d�w� ��f�w���e���N�$�6���!�	�����q���*�l�8�,"B�+"B�k�8��*�r��`   `   �7*���%�+�-�s�>��gS���e�"�r��Hw��r���e��gS�s�>�(�-���%��7*�wD<�ƣX��.x����PU������.x�ģX�wD<�`   `    �9��\.��2�u�>���N�]�\��6d��6d�_�\���N�s�>��2��\.���9�^�V�-"�������E����ƿ��ƿ�E������."��]�V�`   `   U?��\.�)�-�$�6�"�A�x�J�R�M�x�J�"�A�$�6�(�-��\.�U?���e������຿�e�Ol�c�Ol��e��຿������e�`   `    �9���%���!�2�&���-�tj2�rj2���-�4�&���!���%���9���e�)՗�0̿\��-#��5��5��-#�\�0̿*՗���e�`   `   �7*�	��o,�b���S�����S�b��k,�	���7*�^�V�����0̿�E��[6�|7Y��g�{7Y��[6��E�0̿����^�V�`   `   ���?�ԓ������������������ؓ��A����wD<�."���຿\��[6��.g����������.g��[6�\��຿."��yD<�`   `   �����ԾC�ȾS�ž~ržS�žE�Ⱦ��Ծ���q��ƣX������e濩-#�|7Y�����A�������|7Y��-#��e濅���ģX�q��`   `   `����g����/���4����򝾥g��^�������*��.x��E��Ol��5��g����������g��5�Ol��E���.x��*����`   `   P��]O���Mp��k��Mp�]O��%P���x�����l�8������ƿc��5�{7Y��.g�|7Y��5�b���ƿ���l�8������x��`   `   �MX��<��1��1�#�<��MX�?��1ȷ��,"B�PU����ƿOl��-#��[6��[6��-#�Ol���ƿQU��+"B��2ȷ�?��`   `   �;�ņ�l��ņ��;��@�{���K��B!�+"B�����E���e�\��E�\��e濺E�����+"B�E!��K��u���@�`   `   �VؽS���D����Vؽ�k��4�ȹ��K���k�8��.x������຿0̿0̿�຿�����.x�l�8���K��ӹ��4��k�`   `   �����Z������j���� ��4�x��2ȷ������*�ģX�."������*՗�����."��ģX��*�����2ȷ�u���4�� �j���`   `   �&k��&k��ƌ�g����k��@�?���x�����r��wD<�]�V���e���e�^�V�yD<�q������x��?���@��k�j����ƌ�`   `   oM-��<C�Y����(���V��)J��3��3(��Ƨ���\���0�H�B��#I�H�B���0��\�˧��3(���3���)J��V��(��O����<C�`   `   �<C��l�A��cM��� ��+]�����h��h�ɳ�B[�X  �X  �C[�ɳ��g��h������+]��� �\M�A���l��<C�`   `   Y���A��&Խ�l��{@�_�|������*žnD�z��p���Z�o��z��qD��*ž����_�|��{@��l�%ԽA��Y���%�s�`   `   �(��cM��l�78��^l�������-پ����ʈ�������ˈ������-پ������^l�78��l�\M佡(��eN��bN��`   `   �V��� ��{@��^l�`������`$վ(^���
	��>��x��>��
	�(^��]$վ����d���^l��{@��� ��V����0����`   `   �)J��+]�_�|����������Ծ� �����X��������X���� ����Ծ�������c�|��+]��)J��m@�Q�<�S�<��m@�`   `   �3�����������`$վ� ��{�g[�M&��)�M&�g[�}{�� ��c$վ����������3���|��Xэ����Vэ��|��`   `   3(���h���*ž�-پ(^����g[��)��/��/��)�i[���%^���-پ�*ž�h��2(��;�ƾ&�Ѿr�ؾs�ؾ'�Ѿ9�ƾ`   `   Ƨ��h�nD������
	��X�M&��/��Y3��/�M&��X��
	�����lD�h�ȧ��K��dN���!��a&���!�eN�K��`   `   �\�ȳ�z��ʈ��>�����)��/��/��)�����>�ˈ�{��ɳ��\�V�0��O���j�Ș{�Ș{���j��O�V�0�`   `   ��0�B[�p������x����M&��)�M&�����x����o��B[���0�
�Y�xi��eآ�_�����`��eآ�wi��
�Y�`   `   H�B�X  ��Z�����>��X�g[�i[��X��>�����Z�X  �G�B��e|��6��B�ԿW ��{��{�W �B�Կ�6���e|�`   `   �#I�X  �o��ˈ��
	���}{����
	�ˈ�o��X  ��#I�`���&��� �s&�E��#Q�E�s&�� ��&��`��`   `   H�B�C[�z������(^��� ��� ��&^������{��B[�G�B�`��=�ſ���`qE��}��������}�_qE����>�ſ`��`   `   ��0�ɳ�qD辮-پ]$վ��Ծc$վ�-پlD�ɳ���0��e|��&������Q��(��`��@M��`���(���Q�����&���e|�`   `   �\��g��*ž�������������*žh��\�
�Y��6��� �`qE��(���N��+_��+_���N���(��_qE�� ��6���Y�`   `   ˧���h���������d����������h��ȧ��V�0�xi��B�Կs&��}�`��+_��7��+_��`���}�s&�B�Կwi��V�0�`   `   3(�����`�|��^l��^l�d�|����2(��K���O�eآ�W �E����@M��+_��+_��@M�����E�W �eآ��O�J��`   `   �3���+]��{@�78��{@��+]��3��;�ƾdN���j�_���{��#Q����`���N��`������#Q��{�_����j�eN�;�ƾ`   `   �)J��� ��l��l��� ��)J��|��&�Ѿ��!�Ș{�����{�E��}��(���(���}�E��{����Ș{���!�'�Ѿ�|��`   `   �V�]M�&Խ]M��V��m@�Xэ�r�ؾ�a&�Ș{�`��W �s&�_qE��Q�_qE�s&�W �_��Ș{��a&�r�ؾTэ��m@�`   `   �(��A��A���(����Q�<����s�ؾ��!���j�eآ�B�Կ� �������� �B�Կeآ���j���!�r�ؾ���S�<���`   `   O����l�Y���eN���0��S�<�Vэ�'�ѾeN��O�wi���6���&��>�ſ�&���6��wi���O�eN�'�ѾTэ�S�<��0��eN��`   `   �<C��<C�%�s�bN�����m@��|��9�ƾK��V�0�
�Y��e|�`��`���e|��Y�V�0�J��;�ƾ�|���m@���eN��4�s�`   `   ����(�vJj�뿯�f���TD�P���ͯ��c���Z ��>��&S���Z��&S��>�Z �e���ͯ��N����TD�j��뿯�mJj��(�`   `   �(��wL�1����'ǽ�FmF��E��+���0cھ���6��^��^��6���.cھ+����E��GmF���'ǽ3����wL��(�`   `   vJj�1������P�����wP��v�����Oľj�޾��[�����j�޾Rľ����v���wP����P����1���pJj�Y�[�`   `   뿯��'ǽP�����.�7���d������Y��������ξ�Qؾ�Qؾ��ξ�����Y��������d�+�7����R��'ǽ뿯��ऽ�ऽ`   `   f�����.�7���Y�ٹ���n��Γ���F����;b8Ҿ��;�F��Γ���n��ٹ����Y�.�7����h��q ��{��q �`   `   �TD�EmF��wP���d�ٹ�������?�����̾�*վ�*վ��̾@����󩾙��ع����d��wP�FmF��TD��ZF���H���H��ZF�`   `   P����E���v�������n����A��,ξN�پ�0޾Q�پ,ξ>���󩾽n�������v���E��P���!3��=~���S��<~��!3��`   `   ͯ��+�������Y��Γ��?���,ξܾF��E��
ܾ,ξ@���͓���Y�����+���ͯ���ؾR?�������S?��ؾ`   `   c���0cھOľ�����F����̾N�پF��̴�F��N�پ��̾�F������Oľ0cھc����g�X/�oeA��#H�oeA�X/��g�`   `   Z ���j�޾��ξ��;�*վ�0޾E��F�㾿0޾�*վ��;��ξk�޾��Z ��fI�iJw���uG��uG����iJw��fI�`   `   �>��6���Qؾb8Ҿ�*վQ�پ
ܾN�پ�*վe8Ҿ�Qؾ��6��>�P�|��A��)ͿJ쿹���K�)Ϳ�A��P�|�`   `   �&S��^�[����Qؾ��;��̾,ξ,ξ��̾��;�Qؾ[����^��&S�0`����ο��	��*���>���>��*���	���ο0`��`   `   ��Z��^��𾷗ξ�F��@���>��@����F����ξ��^���Z��+���:*���d�ݖ��1��ݖ����d��:*����+��`   `   �&S��6�j�޾����Γ���󩾆�͓������k�޾�6��&S��+�����`�>�����q��O���O���q������`�>�����+��`   `   �>���Rľ�Y���n������n���Y��Oľ���>�0`����`�>����������"��q'��"���������`�>���0`��`   `   Z �.cھ�������ٹ��ع���������0cھZ �P�|���ο�:*���������cm'��lN��lN�cm'����������:*���οQ�|�`   `   e���+����v����d���Y���d��v��+���c����fI��A����	���d�q���"��lN��xe��lN��"�q����d���	��A���fI�`   `   ͯ���E���wP�,�7�.�7��wP��E��ί���g�iJw�)Ϳ�*�ݖ��O����q'��lN��lN��q'�O���ݖ���*�)ͿiJw��g�`   `   N���GmF���������GmF�P����ؾX/���J���>�1��O����"�cm'��"�O���1����>�J���X/��ؾ`   `   �TD��Q��S����TD�!3��R?�oeA�uG��������>�ݖ��q����������q��ݖ����>�����uG��neA�S?�#3��`   `   j���'ǽ����'ǽh���ZF�=~������#H�uG��K��*���d���������������d��*�J�uG���#H����;~���ZF�`   `   뿯�3���1���쿯�q ���H��S�����oeA���)Ϳ��	��:*�`�>�`�>��:*���	�)Ϳ��neA�����S����H�q �`   `   nJj��wL�pJj��ऽ�{����H�<~��S?�X/�iJw��A����ο�������ο�A��iJw�X/�S?�;~����H��{���ऽ`   `   �(��(�Y�[��ऽq ��ZF�!3���ؾ�g��fI�P�|�0`���+���+��0`��Q�|��fI��g��ؾ#3���ZF�q ��ऽ]�[�`   `   �a�`��P-X��C���q ���A�yq���bƾ���'%)��J�5�b�qk�5�b��J�'%)�����bƾzq����A��q ��C��T-X�`��`   `   `��Hi7��,z�Bp��Cm�'u7�Ea|�L����Ӿc�����{x�|x���a�����ӾM��Fa|�%u7�Dm�Dp���,z�Ki7�e��`   `   P-X��,z�lڛ��8˽�����1��e�8������� �žh�־D�ܾe�־ �ž����8����e���1�����8˽nڛ��,z�I-X��^M�`   `   �C��Bp���8˽���>��mZ4��n[�{+��5��uʣ�0׫�1׫�wʣ�5��y+���n[�pZ4�?�����8˽Dp���C��;���:���`   `   �q �Cm����>����%�Ж?��b]��y{����>���I���>�������y{��b]�Ж?���%�>�����Cm��q �I�\��I�`   `   ��A�'u7���1�mZ4�Ж?�TDR�'i���� "��h8��g8���!�����'i�PDR�і?�pZ4���1�%u7���A�V�L��S��S�U�L�`   `   yq��Ea|��e��n[��b]�'i��2z��B拾�+��D拾��2z�'i��b]��n[��e�Ea|�yq�����X慨�T��X慨���`   `   �bƾL��8���{+���y{���������p:��o:�����������y{�y+��7���M���bƾ��较����������`   `   �����Ӿ����5����� "��B拾p:��Ơ��p:��D拾 "�����5��������Ӿ���|�$�lD��;[���c��;[�kD�|�$�`   `   '%)�c��� �žuʣ�>���h8���+��o:��p:���+��g8��?���wʣ��ža���'%)��^��u���N��7���7����N���u���^�`   `   �J���h�־0׫�I���g8��D拾����D拾g8��J���0׫�g�־��	�J�Yo��B���}U����)���}U�B���Yo��`   `   5�b�{x�D�ܾ1׫�>��� "���� "��?���0׫�C�ܾ|x�5�b��~���[��$�WP���k���k�WP���$��[��~��`   `   qk�|x�e�־wʣ��������2z�������wʣ�g�־|x�qk��۶�=`�h�O�-r��yȵ����yȵ�-r��h�O�<`��۶�`   `   5�b��� �ž5���y{�'i�'i��y{�5���ž��5�b��۶�����mk�����=�z/�z/��=�����mk�����۶�`   `   �J�a�������y+���b]�PDR��b]�y+������a���	�J��~��=`��mk��|��P���Y��?r���Y�P��|���mk�=`��~��`   `   '%)���Ӿ8����n[�Ж?�і?��n[�7�����Ӿ'%)�Yo���[�h�O����P�)8r���������)8r�P����h�O��[�Yo��`   `   ���M���e�pZ4���%�pZ4��e�M������^�B�����$�-r���=���Y�����c[��������Y��=�-r����$�A����^�`   `   �bƾFa|���1�@��?����1�Fa|��bƾ|�$��u��}U�WP�yȵ�z/��?r����������?r�z/�yȵ�WP�}U��u��{�$�`   `   zq��&u7���������&u7�yq�����lD��N������k����z/���Y�)8r���Y�z/������k����N��lD����`   `   ��A�Dm��8˽�8˽Cm���A�������;[�7����)���k�yȵ��=�P�P��=�yȵ���k��)�7����;[������`   `   �q �Dp��nڛ�Dp���q �V�L�X慨����c�7�����WP�-r������|�����-r��WP���7�����c���W慨V�L�`   `   �C���,z��,z��C��I��S��T�����;[��N��}U��$�h�O��mk��mk�h�O���$�}U�N���;[����T���S�I�`   `   T-X�Ki7�I-X�;���\���S�X慨��kD��u��B����[�<`����=`��[�A����u��lD���W慨�S�[��;���`   `   `��e���^M�:���I�U�L�������|�$��^�Yo���~���۶��۶��~��Yo���^�{�$���辋��V�L�I�;����^M�`   `   ���_gJ��=�����K�=�����tfƾ#2��,�uBO�K�h�mr�K�h�vBO��,�"2�tfƾ����K�=�����=��ngJ����`   `   ����(��ud�^<����+�� n�~����̾�������"��#����������̾����� n��
+���d<���ud��(����`   `   _gJ��ud�������Zq��I��YJ�����ᚾ���0þFɾ�0þ���ᚾ����YJ��I�]q��������ud�YgJ��KB�`   `   �=��^<������"ʽF ����H1��!S��&s�.���$���$��.���&s��!S��H1���M �"ʽ���d<���=��[G��\G��`   `   �����Zq�F �8�xz��$��9���K�غX��\]�غX���K��9��$�xz��7�F �jq�������] ���] �`   `   K�=�+��I���xz��H��
!�D~-��38�'Y>�$Y>��38�I~-��
!��H�{z����I��
+�M�=�%2N���W���W�"2N�`   `   ����� n��YJ��H1��$��
!���$��1+��0���2��0��1+���$��
!��$��H1��YJ�� n������������9����������`   `   tfƾ~�������!S��9�D~-��1+�n-���.���.�k-��1+�I~-��9��!S��������ufƾ���}�����ߖ�}�����`   `   #2��̾�ᚾ�&s���K��38��0���.�1�.���.��0��38���K��&s��ᚾ�̾!2��*�N��h�ïq��h�N��*�`   `   �,�������.��غX�'Y>���2���.���.���2�$Y>�ܺX�.��볲������,��5h�*���Y���~�¿~�¿Z���*����5h�`   `   uBO�����0þ�$���\]�$Y>��0�l-��0�$Y>��\]��$���0þ���vBO�ނ���:˿T��-B��� �-B�T���:˿ނ��`   `   K�h�"��Fɾ�$��غX��38��1+��1+��38�ܺX��$��Dɾ#��K�h�R���ۈ��^3�ܵd�Ԇ��Ԇ��ܵd��^3�ۈ�S���`   `   mr�#���0þ.����K�I~-���$�I~-���K�.���0þ#��kr�d��Hd��d�����)������)�������d�Hd�d��`   `   K�h�������&s��9��
!��
!��9��&s�볲����K�h�d��q��~��b�������:��:����b�����q��d��`   `   vBO������ᚾ�!S��$��H��$��!S��ᚾ����vBO�R���Hd�~���p����:�.M������.M����:��p��~��Hd�R���`   `   �,��̾����H1�xz�{z��H1�����̾�,�ނ��ۈ��d�b�����:������5���5��������:�b����d�ۈ�߂��`   `   "2������YJ����7����YJ�����!2��5h��:˿�^3��������.M���5��U���5��.M����������^3��:˿�5h�`   `   tfƾ� n��I�N �G ��I�� n�ufƾ�*�*���T��ܵd�)���:������5���5�������:�)��ܵd�T��*����*�`   `   �����
+�]q꽌"ʽkq��
+��������N�Y���-B�Ԇ�������:�.M������.M���:�����Ԇ��-B�Y���N����`   `   K�=�����������M�=����}���h�~�¿�� �Ԇ��)�������:���:����)��Ԇ���� �~�¿�h�}�����`   `   ���d<�����d<�����%2N��������ïq�~�¿-B�ܵd�����b����p��b�������ܵd�-B�~�¿ïq��������%2N�`   `   �=���ud��ud��=���] ���W�8���ߖ��h�Z���T���^3��d���~���d��^3�T��Y����h����7�����W��] �`   `   ngJ��(�YgJ�[G�����W�����}��N�*����:˿ۈ�Hd�q��Hd�ۈ��:˿*���N�}��������W��[G��`   `   �������KB�\G���] �"2N��������*��5h�ނ��S���d��d��S���߂���5h��*�������%2N��] �[G���KB�`   `   JEڼ����,;�1ړ�V��0�3�e��ʽ��� �7^%��|G��,`��>i��,`��|G�7^%��� �ʽ�e��0�3�B��1ړ�#,;�����`   `   ������]O�r-��j�ٽ�	��\��V��ʾ��e��%�o��p���%��e�ʾ��V���\��	�u�ٽ|-���]O������`   `   ,;��]O�тv�=���/z̽���1�A_b�������3s��Q���/s��������A_b��1���3z̽=���тv��]O�,;��5�`   `   1ړ�r-��=����]����ƽ`^�
=�7�-���H�=�^���j���j�B�^���H�/�-�=�q^ｒ�ƽ�]��4���|-��5ړ�>=��@=��`   `   V��j�ٽ/z̽��ƽ��̽�kݽ�)��Wz
��W�Y)"���%�Y)"��W�Wz
��)���kݽĆ̽��ƽHz̽j�ٽH���O������O��`   `   0�3��	���`^��kݽ�\ٽm�߽,��{���������~���7��d�߽x\ٽ�kݽq^����	�2�3��G�=R�=R��G�`   `   e���\��1�
=��)��m�߽�v׽~׽�*ڽK�۽�*ڽ~׽�v׽m�߽�)��
=��1��\�e��m������!J������m��`   `   ʽ��V��A_b�7�-�Wz
�,��~׽VϽ��̽��̽VϽ~׽7��]z
�/�-�=_b��V�� ʽ�"���	������&�`   `   �� �ʾ������H��W�{����*ڽ��̽�[ɽ��̽�*ڽ{����W���H����ʾ��� �i&���I��{c�m��{c��I�i&�`   `   7^%��e����<�^�Y)"����K�۽��̽��̽B�۽���_)"�B�^�����e�8^%�$�a�E��ߩ��������ߩ��E��!�a�`   `   �|G��%�3s����j���%�����*ڽVϽ�*ڽ�����%���j�3s���%��|G��]��8<ƿ����X��~��W������9<ƿ�]��`   `   �,`�o��Q�����j�Y)"�~���~׽~׽{���_)"���j�N���p���,`�3���]���.�<^�M}�M}�<^��.�]��4���`   `   �>i�p��/s��B�^��W�7�뽲v׽7���W�B�^�3s��p���>i�컿�R���]�)P���]�������]��)P����]��R�컿`   `   �,`��%������H�Wz
�d�߽m�߽]z
���H�����%��,`�컿�p��|����$T��2��2�#T�����|��p�컿`   `   �|G��e辷��/�-��)��x\ٽ�)��/�-�����e��|G�3����R��|�!����}2��7u��Z���7u��}2�!����|��R�3���`   `   7^%�ʾ�B_b�=��kݽ�kݽ
=�=_b�ʾ�8^%��]��]����]�����}2�<U���u���u��<U���}2������]�]���]��`   `   �� ��V���1�q^�Ć̽q^��1��V���� �$�a�8<ƿ�.�)P��$T��7u��u��[���u���7u�$T�)P���.�8<ƿ$�a�`   `   ʽ��\�����ƽ��ƽ���\� ʽ�i&�E������<^��]���2��Z���u���u���Z���2��]��<^�����E��j&�`   `   e���	�3z̽�]��Hz̽�	�e��"辁�I�ߩ��X��M}������2��7u�<U���7u��2�����M}�W��ߩ����I�"�`   `   0�3�u�ٽ>���4���j�ٽ2�3�m�����{c����~��M}��]��#T��}2��}2�$T��]��M}�~������{c���k��`   `   B��|-��тv�|-��H�齟G�����	��m����W��<^�)P�����!������)P��<^�W�����m�	�������G�`   `   1ړ��]O��]O�5ړ��O��=R�!J�����{c�ߩ�������.���]��|��|���]��.�����ߩ���{c�	��J��=R��O��`   `   $,;��,;�>=�����=R��������I�E��9<ƿ]���R��p��R�]��8<ƿE����I�������=R����>=��`   `   ���������5�@=���O���G�m��&�i&�!�a��]��4���컿컿3����]��$�a�j&�"�k���G��O��>=���5�`   `   �������&��τ�,ӽQ�"�;�q�,����V�;���3���H�Y�P���H��3�;���V�,���J�q�Q�"�ӽ�τ���&����`   `   ����w��D6�Fk������:�$�C���� ����Ͼ0��:���:��0��Ͼ�������C��:�����Sk���D6��w� ��`   `   �&��D6���U�����y���Y�轠���DC�p�n��ኾ.b��&<��*b���ኾw�n��DC����Y�����������U��D6�~�&���!�`   `   �τ�Fk�������w�����^ý�[�7����$�x 7�bMA�dMA�~ 7���$�.���[�sý���~w������Sk���τ�M���Q���`   `   ,ӽ���y������T���uʩ�Tm����Ͻ�D�r9����r9�D住�Ͻsm��uʩ�0�������������ӽ���Q潊�`   `   Q�"��:�Y��^ýuʩ��>������/��/*��r9��o9��5*���/������>���ʩ�sýN���:�T�"�M6��cA��cA��L6�`   `   ;�q�$�C�����[�Tm�����S��~8��b��b�`��~8�� S�����Ym���[콛��$�C�B�q��ƍ��������������ƍ�`   `   ,�������DC�7����Ͻ�/��~8����i� r^�r^���i�r8���/����Ͻ.���DC����.���Z\Ӿn$��Oj�Nj�m$��_\Ӿ`   `   �V� ���p�n���$��D�/*��b�� r^���S� r^�q��/*���D位�$���n� ����V辩~���6�N�	�V�N���6��~�`   `   ;���Ͼ�ኾx 7�r9�s9��b�r^� r^�V�o9���9�~ 7��ኾ�Ͼ;��[sK�v���C����c���c��D���v���YsK�`   `   �3�0�.b��bMA����o9��`����i�q��o9��׮��bMA�.b��0�3�Od��ޟ���k�����	����k�ߟ��Od��`   `   ��H��:��&<��dMA�r9�5*��~8��s8��/*���9�bMA�$<���:����H�[8��[�޿uS�8y?�\qX�]qX�8y?�tS�[�޿\8��`   `   Y�P��:��*b��~ 7��D��/�� S���/���D�~ 7�.b���:��W�P�3>���Y���>��M���}��Y	���}���M����>��Y�3>��`   `   ��H�0��ኾ��$���Ͻ��������Ͻ��$��ኾ0��H�3>���(�S:W�D-��������������D-��S:W��(�2>��`   `   �3��Ͼw�n�.��sm���>��Ym��.����n��Ͼ�3�[8���Y�S:W�P����q�>��OS�>��q�P���S:W��Y�[8��`   `   :������DC��[�vʩ��ʩ��[��DC� ���;��Od��[�޿��>�D-���q�RES���������RES��q�D-����>�[�޿Od��`   `   �V�������tý1���tý�������V�[sK�ޟ��uS��M������>������M������>������M��uS�ޟ��[sK�`   `   ,����C�Z��������N��$�C�-����~�v����k�8y?��}�����OS����������OS����}��8y?��k�v����~�`   `   J�q��:����~w�������:�B�q�Z\Ӿ��6�C�����\qX�Y	����>�RES�>���Z	��\qX���C�����6�Z\Ӿ`   `   Q�"����������������T�"��ƍ�n$��N��c����	�]qX��}�������q��q������}��\qX���	��c��N�m$���ƍ�`   `   ӽSk����U�Sk��ӽ M6�����Oj�	�V��c����8y?��M��D-��P���D-���M��8y?����c���V�Oj����� M6�`   `   �τ��D6��D6��τ��ὠcA�����Nj�N�D����k�tS���>�S:W�S:W���>�uS��k�C���N�Oj������cA���`   `   ��&��w�~�&�M����Q潞cA�����m$����6�v���ߟ��[�޿�Y��(��Y�[�޿ޟ��v�����6�m$�������cA��Q�M���`   `   ��� ����!�Q������L6��ƍ�_\Ӿ�~�YsK�Od��\8��3>��2>��[8��Od��[sK��~�Z\Ӿ�ƍ� M6���M�����!�`   `   i��������!�Z^a�c��V�*[N�G���zľ�5��y���T'��-��T'�|���5��zľG���<[N�V��b��Z^a��!�����`   `   ����"$ݼ�N�>\��	���뽼,%�t�^�n���ȭ�#�ƾ�Ծ�Ծ$�ƾ�ȭ�o����^��,%����	��^\��N�$ݼ
���`   `   �!��N��N0�<�[�͏��k���D���T!��E�[�e��|�����|�[�e��E��T!��D���k��"͏�<�[��N0��N��!����`   `   Z^a�>\�<�[�ǣg��@��{I���Ժ��\�������������������\ཙԺ��I���@����g�#�[�_\�c^a���e���e�`   `   c���	��͏��@����x�â~����dt������E����ζ�E�������dt��:���â~�n�x��@��?͏��	���b��������ƽ����`   `   V����k��{I��â~�3�^�Q��8P�&�T���X���X�3�T��8P��Q��^��~��I���k����V��(�V6'�S6'��(�`   `   *[N��,%��D���Ժ����Q�mj)�d������	����d��lj)�Q�����Ժ��D���,%�3[N��os�f����i��k����os�`   `   G���t�^��T!��\�dt���8P�e����"
˼=
˼��I���8P�tt���\��T!���^�H����)���о+�߾'�߾�о�)��`   `   zľn���E��������&�T����"
˼ݳ��"
˼܎�&�T�|������%�E�n��zľrD�����-� 4��-���rD��`   `   �5���ȭ�Z�e���E�����X��	�=
˼"
˼�	���X�U������T�e��ȭ��5���3*���X�(s��j��k��*s����X��3*�`   `   y��#�ƾ�|�����ζ���X������܎���X��ζ�����|�#�ƾ{��!{V�2���L�����ѿ)ܿ��ѿL���4���!{V�`   `   �T'��Ծ������E���4�T�e��I��&�T�U����������Ծ�T'�|�Q/��S^�d��n&�o&�e��Q^�P/��|�`   `   �-��Ծ�|���������8P�mj)��8P�|�������|��Ծ߿-������Ͽ(L�*�E���n��|���n�+�E�(L��Ͽ����`   `   �T'�$�ƾZ�e����dt���Q�Q�tt�����T�e�#�ƾ�T'�����}2ٿ�h%��Yn��;��+͹�+͹��;���Yn��h%�}2ٿ����`   `   |���ȭ��E��\�:����^�����\�%�E��ȭ�{��|��Ͽ�h%�b�~�<����l���5��l��<���a�~��h%��Ͽ|�`   `   �5��o���T!��Ժ�â~��~��Ժ��T!�n���5��!{V�Q/��(L��Yn�<���-�*u$�*u$�-�<����Yn�(L�P/��"{V�`   `   zľ��^��D���I��n�x��I���D����^�zľ�3*�2���S^�*�E��;���l��*u$���6�*u$��l���;��*�E�S^�2����3*�`   `   G����,%��k���@���@���k���,%�H���rD����X�L���d����n�+͹��5�*u$�*u$��5�+͹���n�e��L�����X�tD��`   `   <[N���"͏���g�?͏���3[N��)����(s����ѿn&��|�+͹��l��-��l��+͹��|�n&���ѿ(s�����)��`   `   V��	��<�[�#�[��	��V��os��о�-�j��)ܿo&���n��;��<���<����;����n�n&�)ܿk���-��о�os�`   `   �b��_\��N0�_\��b���(�f���+�߾ 4�k����ѿe��+�E��Yn�a�~��Yn�*�E�e����ѿk�� 4�+�߾k����(�`   `   Z^a��N��N�c^a�����V6'��i��'�߾�-�*s��L���Q^�(L��h%��h%�(L�S^�L���(s���-�+�߾�i��S6'�����`   `   �!�$ݼ�!���e���ƽS6'�k����о����X�4���P/���Ͽ}2ٿ�ϿP/��2�����X����оk���S6'���ƽ��e�`   `   ����
��������e������(��os��)��rD���3*�!{V�|���������|�"{V��3*�tD���)���os��(�������e�Ǔ�`   `   �,W�������Ӽ�D1�r"��\�߽�%�
�h�����~�ľ��龟�r�������~�ľ����
�h��%�\�߽O"���D1�۶Ӽ����`   `   ����ޚ��q漓L+���������U�|�0��Ob�����E��eʦ�iʦ�F�������Ob���0��U�����­��L+��p�Ú������`   `   ��Ӽq�ï���(�>S^�Ɣ�i�Ľ���aq�y�3���D��K���D�y�3�iq����]�ĽƔ�NS^���(����q演�ӼiMμ`   `   �D1��L+���(�l�/���C�8Eg�u>���\ŽG\ܽMA�PA�V\ܽ\Ž�悔f>��oEg���C�9�/���(��L+��D1���5���5�`   `   r"�����>S^���C�iO5���4���@���T�E�i��z�����z��i���T��@���4�O5���C��S^����\"�����ja�����`   `   \�߽����Ɣ�8Eg���4�5T�
m�����i�������������ъ���l�T���4�oEg�Ɣ�����`�߽����Y��Y�m���`   `   �%��U�i�Ľu>����@�
m�J���������l�:*`���l�����J���
m���@�u>��[�Ľ�U��%�j�C� Y�!�`�Y�j�C�`   `   
�h�|�0����𨽀�T���������@���㻻任$������ъ����T��悔�����0��h�`Ǐ�2ե�f=��b=��0ե�fǏ�`   `   �����Ob�aq�\ŽE�i�i����l��㻻/ME��㻻��l�i���i�\Žsq��Ob�����"�Ⱦ�����v�������"�Ⱦ`   `   ~�ľ����y�3�G\ܽ�z�����:*`�任�㻻�)`������z�V\ܽs�3������ľL����'�{�D���U���U�~�D���'�H��`   `   ���E����D�MA齖��������l�$����l��������MA齹�D�E�����`r%���[�^���n��,����n��^����[�`r%�`   `   ��eʦ��K�PA��z������������i���z�MA��K�iʦ���b�@�.���l�����տ�m쿐m���տk���-���e�@�`   `   r��iʦ���D�V\ܽ�i�ъ��J���ъ���i�V\ܽ��D�iʦ�p���dP�U����Կ9^	�O�!��[+�O�!�9^	���ԿU���dP�`   `   ��F��y�3�\Ž��T��l�
m���T�\Žs�3�E�����dP�>2��z��bn!� QL��h��h� QL�bn!�|��>2���dP�`   `   �������iq��悔�@�T���@��悔sq��������b�@�U��z��¿*���g�l��o_��l����g���*�z��U��b�@�`   `   ~�ľ�Ob����f>����4���4�u>������Ob��ľ`r%�.�����Կbn!���g��Q������ߝ���Q����g�bn!���Կ-���ar%�`   `   ������0�]�ĽoEg�O5�oEg�[�Ľ��0�����L����[�l���9^	� QL�l��������������l�� QL�9^	�l�����[�L��`   `   
�h��U�Ɣ���C���C�Ɣ��U��h�"�Ⱦ��'�^����տO�!��h�o_��ߝ������p_���h�O�!���տ^����'�$�Ⱦ`   `   �%�����NS^�9�/��S^������%�`Ǐ����{�D��n���m��[+��h�l���Q��l���h��[+��m��n��{�D����`Ǐ�`   `   \�߽­���(���(����`�߽j�C�2ե�����U�,����m�O�!� QL���g���g� QL�O�!��m�,�����U���0ե�b�C�`   `   O"���L+�����L+�\"������Y�f=��v����U��n����տ9^	�bn!���*�bn!�9^	���տ�n����U�s��f=��
Y����`   `   �D1��p�q漢D1�����Y�!�`�b=����~�D�^��k�����Կ|��z�꿷�Կl���^��{�D���f=���`��Y���`   `   ۶ӼÚ����Ӽ��5�ja���Y�Y�0ե���񾐸'���[�.���U��>2��U��.�����[���'����0ե�
Y��Y�_a����5�`   `   ��������iMμ��5����m���j�C�fǏ�"�ȾH��`r%�e�@��dP��dP�b�@�ar%�L��$�Ⱦ`Ǐ�b�C��������5�4Mμ`   `   
�޻�������y���W�S���.�����-�5g�^�)��{���@ľ{����)��^#g���-�X������S�y���׍�����`   `   ���rH�������>9��e����½f:��'�VJ���e��9u��9u���e�VJ���'�t:���½�e��b9�A��ޭ���qH���`   `   ����������������U�f����ʷ���ὙK����������K�����ʷ�Z����U� ����}�����������w��`   `   z�����（�鼾�������LB��l������~���夽�夽�~�������l��KB�)��A��T��R��A�＋����_��_�`   `   W�S�?9�������K��p&�����Q��=��w�#�=��#�����'��K�������_�?9�)�S��g�vn��g�`   `   ���e���U����K�缭.��OW���dx��	p���o�x�o��	p�[ex�W��K.�����)��ϓU��e���������˽�˽����`   `   .�����½g���LB�p&��OW�����jMd�!�m�����m�jMd����OW���&��LB�X�����½E���qF�E_#�C!)�R_#�qF�`   `   ��-�f:��ʷ��l�����dx�kMd��6`;�;��;@7`;uKd�[ex�����l��ʷ�t:���-���V�l�w�B߄�>߄�h�w���V�`   `   5g��'���Ὃ���Q���	p�%�m��;J�<�;��m��	p�����������'�%g�aw�����`�ƾM:ξ`�ƾ~��aw��`   `   ^VJ��K��~��=����o�����;�;E��y�o�`���~���K�VJ�_�¾���ډ�������݉����¾`   `   �)����e�����夽x�#�y�o���m�?7`;��m�y�o�[�#��夽�����e��)��V"����"?��5X��na��5X��"?����V"�`   `   {����9u����夽=���	p�lMd�wKd��	p�`���夽ۂ��9u�|���
�D>=�:�r��k�����������k��6�r�C>=�
�`   `   @ľ�9u�����~��#��\ex����\ex����~������9u�;ľ$��@�T�ۑ���@��п��ڿп�@��ۑ��>�T�$��`   `   {�����e��K��������W��OW����������K���e�|���$��6�]�����xjϿڡ��������١��zjϿ����5�]�"��`   `   �)��VJ���Ὃl�'��L.���&���l����VJ��)��
�@�T�����_�ٿ���F4&�i0�H4&����\�ٿ����C�T�
�`   `   ^��'��ʷ��KB�K�缒��LB��ʷ��'�_V"�D>=�ۑ��xjϿ���0�s`F�s`F�0����zjϿڑ��C>=�W"�`   `   #g�t:�Z���)�����)��W���t:�%g��¾��:�r��@��ڡ��F4&�s`F�\S�s`F�F4&�ڡ���@��:�r�����¾`   `   ��-���½�U�A����ϓU���½��-�aw������"?��k��п���i0�s`F�s`F�j0����п�k���"?����cw��`   `   X����e�� �T��_��e��D�����V����ډ��5X�������ڿ���H4&�0�F4&������ڿ�����5X�ډ������V�`   `   ��b9����R��>9���pF�l�w�`�ƾ����na�����п١��������ڡ��п�����na����b�ƾh�w�iF�`   `   �S�A��}���A��)�S�����E_#�B߄�M:ξ����5X��k���@��zjϿ\�ٿzjϿ�@���k���5X����G:ξB߄�Q_#�����`   `   y���ޭ����������g��˽C!)�=߄�`�ƾ݉��"?�6�r�ۑ����������ڑ��:�r��"?�ډ�b�ƾB߄�;!)��˽�g�`   `   ׍���qH������_�vn��˽R_#�h�w�~��������C>=�>�T�6�]�C�T�C>=���������h�w�Q_#��˽bn��_�`   `   ������w���_��g�����pF���V�aw���¾V"�
�$��"��
�W"ﾡ¾cw����V�iF������g��_��w��`   `   �����'��@�A ��aX
�q.c�u^��z�0	 ���G�f�j�1���a݅�1���p�j���G�	 �z�^��q.c�X
�A ��*A��'�`   `   �'�Bo���y������{뼬�6��F�����j��12�;���Y(��Y(�<��%2�r������F��x�6�*|�����Gy��n��(�`   `   �@��y���@���������F��:�K�t�\���3R���½yɽ�½3R��l���K�t���:�F�ǀ��������@��y��@�����`   `   A ������������������(���s�By��/�[=F��4S��4S�x=F��/�y��s뼗��𐙼$����������R ���i���i��`   `   aX
��{뼦��������K��c[m���v�����ɛ�5��G��5�]ɛ������v�c[m�K������C����{�4X
�C��CJ�C��`   `   q.c���6�F�(��c[m��=��y����E����#K��J����k�E��x��=��[m����+�x�6�y.c��+���㌽�㌽�+��`   `   u^���F���:��s뼐�v��y���;\O�;�~<��<�~<]O�;��;�y����v��s���:��F���^���Dͽ!n佭��;n��Dͽ`   `   z����K�t�Cy������E�\O�;D<�o<�o<D<XP�;l�E���y�1�t����z�2��ƣ,�:M9�1M9�ã,�?��`   `   0	 �j��]����/��ɛ�����~<�o<kQ�<�o<-~<���8ɛ��/�����j�� 	 �ĤM�_�u��ሾ�፾�ሾV�u�ĤM�`   `   ��G�12�3R��[=F�6�%K���<�o<�o<C�<�J�|�x=F�&R��%2���G�~1��'}�������Dξ�Dξ����%}��w1��`   `   f�j�;���½�4S��G���J��~<D<-~<�J��G���4S��½;��p�j�τ���1ҾP����D�����D�P����1Ҿτ��`   `   1����Y(�yɽ�4S�6����[O�;WP�;���|��4S�lɽ�Y(�2���$��g���\�0G9���H���H�3G9�X�e���$��`   `   a݅��Y(��½x=F�]ɛ�m�E���;m�E�8ɛ�x=F��½�Y(�\݅��lǾg���	8�,�a��Y���	���Y��-�a��	8�e���lǾ`   `   1���<��3R���/�����x���y�����/�&R��;��2����lǾ��e G�����w�����������w�����h G����lǾ`   `   p�j�%2�l���y���v�=���v�y�����%2�p�j�$��g��e G�Ce�������߿� Xɿ�߿�����@e��e G�i��$��`   `   ��G�r��K�t��s�c[m��[m��s�1�t�j�潰�G�τ��g����	8���������<ɿ�޿�޿�<ɿ��������	8�e���Є��`   `   	 ������:����K�������:���� 	 �~1���1Ҿ\�,�a��w���߿��޿�u鿊޿�߿��w��+�a�\��1Ҿ~1��`   `   z��F��F�𐙼����+��F��z�ĤM�'}��P���0G9��Y������ Xɿ�޿�޿Xɿ�����Y��3G9�Q���%}��ȤM�`   `   �^��x�6�ǀ��$���C���x�6��^��2��_�u������D���H��	�������߿��<ɿ�߿������	����H��D�����_�u�2��`   `   q.c�*|뼴�������{�y.c��Dͽƣ,��ሾ�Dξ�����H��Y���w�����������w���Y����H�����Dξ�ሾ£,��Dͽ`   `   X
�������@�����4X
��+��!n�:M9��፾�Dξ�D�3G9�-�a����@e�����+�a�3G9��D��Dξ�፾:M9�8n佫+��`   `   A ��Gy��y�Q ��C���㌽���1M9��ሾ����P���X��	8�h G�e G��	8�\�Q��������ሾ:M9���콄㌽f��`   `   *A��n���@��i��CJ��㌽;n�£,�V�u�%}���1Ҿe���e����i��e����1Ҿ%}��_�u�£,�8n佄㌽/J��i��`   `   �'�(������i��C���+���Dͽ?��ĤM�w1��τ��$���lǾ�lǾ$��Є��~1��ȤM�2���Dͽ�+��f���i������`   `   �u�;0̑;pK�9�
㻥��wO�ŠT�����D`̽����H>%�Ϊ*�H>%�#����"`̽�����T�wO����
㻣7�90̑;`   `   0̑;��<;Z����Ż>�g���̼�����]��N��x���ǽv&ս�&ս�ǽx���N����]�d����̼Ŷg���Ż��s�<;�ˑ;`   `   eK�9^�����nY��!$&�yd����ͼ�l�o^4��V��m�=u��m��V��^4��l���ͼyd��[$&�nY��(��_���H�9�:`   `   �
㻐�ŻoY��������׻�����S��m���Ӵ�]Ӽ�����㼑ӼԴ�em��k�S�x��Н׻x����X����Ż9�3�������`   `   ���>�g�!$&���׻�΄�"�:�kR>��z�h���@Ȼf1ջ�@Ȼ�f���z�W>�"�:�̄���׻J%&�>�g�P��^^��"��^^��`   `   wO���̼yd�����#�:��J�:lך;[��;��;��;��;���;���;aؚ;P�:A�:�y��Fd����̼O�7���,���,��6�`   `   ŠT������ͼ��S�mR>�kך;��$</\<νy<Lx�<�y</\<��$<kך;S>���S���ͼ����T��ǁ�?���9[��X����ǁ�`   `   ������]��l��m���z�Z��;/\<�j�<
�<�	�<�j�<�\<���;5�z�fm���l���]�����5��]�޽��ｕ��V�޽+5��`   `   D`̽�N��o^4��Ӵ�h����;νy<
�<���<
�<D�y<��;2f���Ӵ��^4��N��&`̽9I��s��h0�'�6��h0��s�9I�`   `   ���x���V�]Ӽ�@Ȼ��;Lx�<�	�<
�<�x�<��;�AȻ�Ӽ�V�x�����i�*���S�;t�����Gt���S�\�*�`   `   ��ǽ�m����h1ջ��;�y<�j�<C�y<��;y0ջ��㼾m��ǽ"��2O����W@������1�����W@�����2O�`   `   H>%�v&ս=u���㼬@Ȼ���;/\<�\<��;�AȻ����<u��&սJ>%�^l��0����þE�⾧p���p��I�⾺�þ�0��il�`   `   Ϊ*��&ս�m��Ӽ�f�����;��$<���;2f���Ӽ�m��&սƪ*�U*|������I�����������J���ᾒ��U*|�`   `   H>%��ǽ�V�Դ��z�`ؚ;kך;5�z��Ӵ��V��ǽJ>%�U*|�������D����1���@���@���1�F�������O*|�`   `   #�x���^4�fm��W>�P�:S>�fm���^4�x��"�^l�������ݷ��T@�څY���b���Y��T@�ط������^l�`   `   ����N���l�k�S�$�:�A�:���S��l��N������2O��0����D���T@�#�b���v���v� �b��T@�F��ᾁ0���2O�`   `   "`̽��]���ͼy��̄�x����ͼ��]�&`̽i�*������þI����1�څY���v�)�����v�څY���1�I����þ���i�*�`   `   ����d��yd��Н׻��׻Fd���������9I���S�W@��D�⾠����@���b���v���v���b���@����I��X@����S�=I�`   `   �T���̼[$&�x���J%&���̼�T�5���s�;t�����p�������@���Y� �b�څY���@�����p��
���;t��s�5��`   `   wO�Ŷg�nY���X��>�g�O��ǁ�]�޽�h0����1���p�������1��T@��T@���1�����p���1�����h0�V�޽�ǁ�`   `   ����Ż(����ŻP��7�?������&�6������I��J��F��ط�F��I��I��
������6����U���7�`   `   �
����Z��7�^^����,�9[����ｬh0�Gt�W@����þ�ᾌ�񾆭����þX@��;t��h0����*[����,��^��`   `   �7�9s�<;�H�91���"����,�W���V�޽�s���S����0������������0�������S��s�V�޽U�����,����2���`   `   0̑;�ˑ;�:����^^���6��ǁ�+5��9I�\�*��2O�il�U*|�O*|�^l��2O�i�*�=I�5���ǁ�7��^��2���\�:`   `   �A6<,�'<�c�;��);<�����k�2lڼ@)(��h�����l�����z7ǽ����l������h�@)(��lڼ��k�L�����);�b�;,�'<`   `   ,�'<1z<t�;��V;3���b����V��'��ȇA���_���o�	�o���_���A�8�����}��	b�/����V;�t�;`z<
�'<`   `   �c�;t�;7S�;(u~;քa:~Z������m�	ݧ�*Ҽ�������_��*Ҽ4ݧ���m�{��Z��a:(u~;gS�;
t�;�c�;4�;`   `   ��);��V;'u~;��;Y;e;{;��n�F@F��Y�����-��5��*��tZ���=F��wn�-x;\9e;f�;�v~;��V;C�);�a;a;`   `   >���6��΄a:W;e;��;s�;���;���;���;UO�;-�;UO�;߹�;���;���;s�;,!�;X;e;ta:6��	��� �һ�� �һ`   `   ��k��b��Z�{;s�;Ko"<��G<�]<��h<km<km<��h<��]<(�G<�o"<
r�;+x;�Z�
b���k�޾��cH��LH������`   `   3lڼ�������n����;��G<xx�<I�<��<͍�<��<I�<jx�<��G<���;ߔn�i�����wlڼlj��o!�o�(��o!�lj�`   `   @)(�V�Ἤ�m�I@F����;�]<I�<h�<�u�<�u�<!h�<��<��]<���;�=F�K�m����I)(��[��7��z���k����7���[�`   `   �h�(��	ݧ��Y�����;��h<��<�u�<(��<�u�<Y�<��h<X��;�Y���ݧ�'���h��/��s꺽�/ѽ�ٽ�/ѽc꺽�/��`   `   ���ȇA�*Ҽ���TO�;km<͍�<�u�<�u�<��<km<VN�;+���Ҽ��A����b�ȽΏ��s���ʘ�~��ɏ��K�Ƚ`   `   �l����_����.��
-�;km<��<!h�<Y�<km<�-�;-�����_��l��%����%�;���P��_X���P�%�;���%��`   `   �����o�����6��TO�;��h<I�<��<��h<VN�;-������	�o����� �%�8�M�d�Ѳ��,o��2o��Բ��A�d�"�8��`   `   z7ǽ	�o�`��+��޹�;��]<jx�<��]<X��;+�����	�o�k7ǽrZ���K��}��.�)���T+��)���/򛾌}����K�rZ�`   `   �����_�*ҼvZ�����;(�G<��G<���;�Y���Ҽ��_����rZ�6�R����1ᬾ��Ǿ�8׾�8׾{�Ǿ4ᬾ���3�R�mZ�`   `   �l����A�4ݧ��=F����;�o"<���;�=F��ݧ���A��l��� ���K����|���r�־l�u9��w�r�־s��������K�� �`   `   ���8����m��wn�s�;
r�;֔n�K�m�'�����%��%�8��}��1ᬾr�־$
��'I�$I�
��v�־4ᬾ�}��"�8�&��`   `   �h����{��+x;,!�;,x;h����Ἴh�b�Ƚ��M�d�-򛾁�Ǿl�&I�{�&I�l��Ǿ,�M�d���b�Ƚ`   `   @)(�}���Z�\9e;X;e;�Z����H)(��/��Ώ��%�;�в��)����8׾u9��$I�&I�z9���8׾&���Բ��&�;�ȏ���/��`   `   �lڼ	b��a:f�;ta:	b�wlڼ�[�s꺽s����P�,o��T+���8׾w�
��l�8׾\+��,o����P�s��p꺽�[�`   `   ��k�0��(u~;�v~;3����k�lj��7���/ѽ��_X�2o��)���{�Ǿr�־v�־��Ǿ&���,o���_X�ʘ��/ѽ�7��Oj�`   `   M�����V;gS�;��V;���ݾ���o!�y����ٽʘ���P�Բ��/�4ᬾs���4ᬾ,�Բ����P�ʘ��ٽz����o!�ݾ��`   `   ��);�t�;t�;E�);��һcH��o�(�j����/ѽ~��%�;�A�d��}���������}��M�d�&�;�s���/ѽz���R�(�LH����һ`   `   �b�;`z<�c�;�a;��LH���o!��7��c꺽ȏ����"�8���K�3�R���K�"�8���ȏ��p꺽�7���o!�LH��E軾a;`   `   ,�'<
�'<5�;a;��һ����lj��[��/��K�Ƚ%���rZ�mZ�� �&��b�Ƚ�/���[�Oj�ݾ����һ�a;��;`   `   M�}<ӷt<-7X<�K&<���;|�{���1ㅼ�UѼ�R� l,��jA�~�H��jA�?l,��R�:UѼ1ㅼh��������;�K&<�6X<ӷt<`   `   ӷt<I+j<��S<�.<>��;T�Q;���{ ���c��Y���{¼��ռ��ռ�{¼�Y����c��{ ������Q;X��;�.<ޘS<k+j<��t<`   `   -7X<��S<2�I<�S7<^�<Fh�;���;�U�9��G��Oǻ�c��T��c��Oǻ��G��U�9��;Eh�;E�<�S7<;�I<��S<-7X<��Y<`   `   �K&<�.<�S7<)O<<#:<��.<�<�9<���;���;���;���;��;D��;f:<��<:�.<�":<�O<<$T7<�.<`K&<0 !< !<`   `   ���;=��;^�<#:<�}R<�wa<�+g<��e<��a<�>]<�[<�>]<�a<��e<�*g<�wa<�~R<#:<y�<=��; ��;��;�w�;��;`   `   ��Q�Q;Dh�;��.<�wa<�<׀�<3��<�v�<�m�<�m�<�v�<��<��<S�<Zwa<:�.<�h�;��Q;���F�����U�����F�`   `   ~���������;�<�+g<׀�<I7�<M}�<�i�<L�<�i�<M}�<77�<׀�<�+g<�<4��;���R���a�N�@ ������ ��a�N�`   `   2ㅼ{ ��U�9�9<��e<3��<M}�<2��<�<`�<3��<�}�<��<6�e<e:<�`�9�{ �Cㅼ"eżK ��yW�`W�: ��heż`   `   �UѼ��c���G����;��a<�v�<�i�<�</��<�<bi�<�v�<E�a<���;��G���c�JUѼu#��>�4Y�?�b�4Y���>�u#�`   `   �R��Y���Oǻ���;�>]<�m�<L�<`�<�<��<�m�<�>]<��;Oǻ�Y���R���L�����l���ئ�٦��l�� �����L�`   `   !l,��{¼�c����;�[<�m�<�i�<3��<bi�<�m�<t�[<���;�c��{¼7l,�	I~������+ʽ^���@���+ʽ����	I~�`   `   �jA���ռ�T����;�>]<�v�<M}�<�}�<�v�<�>]<���;6T���ռ�jA�4��ƽ�����D��������D�����ƽ"4��`   `   �H���ռ�c���;�a<��<77�<��<E�a<��;�c���ռe�H�������ڽ{����'���:�6/A���:���'�{����ڽ����`   `   �jA��{¼�OǻC��;��e<��<׀�<6�e<���;Oǻ�{¼�jA������:�T2��X9�_>U���d���d�U>U��X9�[2��:�y���`   `   ?l,��Y����G�e:<�*g<S�<�+g<e:<��G��Y��7l,�4����ڽT2��?��d��t}�G��u}��d�q�?�T2���ڽ4��`   `   �R���c��U�9��<�wa<Ywa<�<�`�9��c��R�	I~�ƽ{���X9��d��(�����������(���d��X9�w��ƽ	I~�`   `   ;UѼ�{ ���;:�.<�~R<:�.<4��;�{ �IUѼ��L�����������'�_>U��t}������������t}�_>U�~�'�����������L�`   `   1ㅼ���Eh�;�":<#:<�h�;���Bㅼu#�����+ʽ�D���:���d�G����������G����d���:��D��+ʽ ����#�`   `   h�����Q;E�<�O<<y�<��Q;P���!eż�>��l��^�὿��6/A���d�u}��(���t}���d�C/A����Q�Ὦl���>�!eż`   `   ��X��;�S7<$T7<>��;��`�N�J ��4Y��ئ�������:�U>U��d��d�_>U���:�����٦�4Y�9 ����N�`   `   ���;�.<;�I<�.<��;�F�@ ��xW�?�b�٦�@�ὰD���'��X9�q�?��X9�~�'��D�Q��٦��b�xW�� ���F�`   `   �K&<ޘS<��S<aK&<���;�������`W�4Y��l���+ʽ����{��[2�S2�w�������+ʽ�l��4Y�xW�̅��S������;`   `   �6X<k+j<-7X<1 !<�w�;R���� ��9 ����>� �������ƽ��ڽ�:���ڽƽ���� ����>�9 ��� ��S����x�;0 !<`   `   ӷt<��t<��Y< !<���;��F�`�N�geżu#���L�	I~�"4������y���4��	I~���L��#�!eż��N��F����;0 !<�Y<`   `   ���<S�<Տ<Qz�<��X<�l!<}Y�;2vk:�t��\,���X�E7��49��E7����X�\,��s��0vk:�W�;�l!<u�X<Qz�<�ԏ<S�<`   `   S�<��<�ߎ<E��<̈l<}lF<y�<,��;��0;Fy���C1��䂻K傻cC1��m����0;J��;չ<�lF<h�l<!��<�ߎ<��<B�<`   `   Տ<�ߎ<���<G}�<ג�<��n<6JT<��5<\�<��;&��;C��;v��;��;;�<��5<JJT<��n<Ԓ�<F}�<���<�ߎ<%Տ<S�<`   `   Qz�<E��<F}�<�y�<&�<�ˊ<�{�<�N�<P=s<� h<<�a<C�a<~ h<=s<�N�<�{�<�ˊ<�~�<�y�<n}�<!��<@z�<�*<�*<`   `   ��X<ˈl<ג�<&�<;p�<%��<ҽ�<ʚ�<�,�<,y�<")�<,y�<�,�<ʚ�<v��<%��<�p�<&�<{��<ˈl<3�X<��K<!G<��K<`   `   �l!<|lF<��n<�ˊ<%��<o��<`�<R��<��<�!�<�!�<�<;��<��<���<�<�ˊ<��n<�lF<�l!<W<��;:��;�<`   `   {Y�;x�<5JT<�{�<ҽ�<`�<��<|��<���<���<���<|��<��<`�<ֽ�<�{�<XJT<x�<�X�;�/;@�/:�[�{�/:�/;`   `   vk:)��;��5<�N�<ʚ�<R��<|��<��<*�<�<��<���<;��<���<�N�<F�5<H��;�sk:k�u�P�x;�1;�'��u�`   `   u����0;[�<P=s<�,�<��<���<*�<S��<*�<p��<��<�,�<P=s<��<��0;�s���x1��z��*������*��az���x1�`   `   ^,�my����;� h<,y�<�!�<���<�<*�<ԯ�<�!�<�x�<} h<A�;�m���,�6����ռ�M�o����M���ռ����`   `   ��X��C1�$��;;�a<!)�<�!�<���<��<p��<�!�<W)�<;�a<���;�C1���X���ȼ�0��7�СP�ɦY���P��7��0���ȼ`   `   E7���䂻A��;B�a<,y�<�<|��<���<��<�x�<;�a<���;M傻V7����|y1���e�߆��ᑽ�ᑽ߆�v�e�wy1���`   `   49��M傻u��;} h<�,�<:��<��<:��<�,�<} h<���;M傻9��)��`+G�u���c�2)��q���2)��h�u���N+G�)��`   `   E7��fC1���;=s<ʚ�<��<`�<���<P=s<A�;�C1�V7��)����N��m��]���_�ν\e޽Oe޽Q�νf����m����N���`   `   ��X��m��;�<�N�<v��<���<ֽ�<�N�<��<�m����X���`+G��m��%丽׈ݽ���H|�����׈ݽ丽�m��q+G���`   `   ],���0;��5<�{�<%��<�<�{�<G�5<��0;,���ȼ{y1�u���]���׈ݽ--��p��i�� -���ݽf���o���vy1���ȼ`   `   �s��I��;JJT<�ˊ<�p�<�ˊ<XJT<I��;�s��5����0���e�c�_�ν���p��{��p�����_�ν`򠽒�e��0�5���`   `   )vk:չ<��n<�~�<&�<��n<x�<tk:�x1��ռ�7�߆�2)��\e޽H|��i��p��S|��Oe޽,)��߆��7���ռ�x1�`   `   �W�;�lF<Ԓ�<�y�<{��<�lF<�X�;g�u��z���M�ϡP��ᑽq���Oe޽��� -�����Oe޽�����ᑽ��P��M�xz��h�u�`   `   �l!<h�l<F}�<n}�<ˈl<�l!<�/;M�*��o�ȦY��ᑽ2)��Q�ν׈ݽ�ݽ_�ν,)���ᑽƦY���:*��%�v�/;`   `   u�X<!��<���<!��<4�X<X<R�/:w;���������P�߆�h�f���丽f���`�߆���P���Q���w;�?�/:W<`   `   Qz�<�ߎ<�ߎ<@z�< �K<��;|Z�/;�*���M��7�v�e�t����m���m��o�����e��7��M�9*��w;�E��<��;��K<`   `   �ԏ<��<%Տ<�*<"G<<��;��/:$�`z����ռ�0�vy1�N+G���N�q+G�vy1��0���ռxz��$�A�/:<��;qG<�*<`   `   S�<B�<S�<�*< �K<�<�/;�u��x1�������ȼ��)�������ȼ5����x1�f�u�w�/;X<��K<�*<z�<`   `   Vc�<)��<��<�k�<�ח<��<>�q<�J<� <2��;�;s�};��];s�};��;2��;( <�J<��q<��<�ח<�k�<���<)��<`   `   )��<阬<j��<-�<�d�<]m�<S1�<��z<t�_<P�F<��3<�8)<�8)<ȼ3<��F<@�_<\�z<y1�<m�<�d�<�<���<혬<��<`   `   ��<j��<�Y�<[Q�<^�<��<�M�<7Y�<�<X}�<��<GH�<��<X}�<��<7Y�<�M�<��<d�<[Q�<�Y�<j��<(��<���<`   `   �k�<-�<[Q�<�g�<���<�8�<�U�<3�<�y�<5�<C��<J��<(�<�y�<#3�<�U�<k8�<\��<
h�<{Q�<�<�k�<���<���<`   `   �ח<�d�<]�<���<e�<��<��<��<��<!�<,�<!�<��<��<s�<��<��<���<�<�d�<�ח<�v�<��<�v�<`   `   ��<\m�<��<�8�<��<�{�<���<L��<	��<���<y��<��<>��<���<�{�<��<k8�<��<m�<��<�!�<Ȱx<ΰx<�!�<`   `   =�q<S1�<�M�<�U�<��<���<�y�<�u�<L��<��<m��<�u�<ry�<���<��<�U�<�M�<S1�<�q<XQT<K�@<M�9<�@<XQT<`   `   �J<��z<6Y�<3�<��<K��<�u�<F�<>��<$��<F�<�u�<>��<ܒ�<#3�<WY�<[�z<yJ<�i<Q�;E2�;�2�;Q�;�i<`   `   � <s�_<�<�y�<��<	��<L��<>��<D��<>��<-��<	��<��<�y�<��<s�_< <���;�B;��o:g`F9��o:�B;���;`   `   0��;O�F<X}�<5�<!�<��<��<$��<>��<��<y��<� �<(�<x}�<��F<��;mr ;��ʫ����٣滑ʫ�����s ;`   `   �;��3<��<C��<,�<x��<l��<F�<-��<y��<[�<C��<��<��3<��;��Q���׻�x;�ؕp�<���g�p��x;�Y�׻��Q�`   `   n�};�8)<FH�<J��<!�<��<�u�<�u�<	��<� �<C��<gH�<�8)<�};��U��+�%�������ʼ<�ʼ��� ����+�|�U�`   `   ��];�8)<��<(�<��<>��<ry�<>��<��<(�<��<�8)<��];u���OzV�ف���R��������S�ف��zV�u���`   `   o�};ȼ3<X}�<�y�<��<���<���<ܒ�<�y�<y}�<��3<�};t���Dxe�����` �F}/�5}/�` ���+��=xe�@���`   `   ��;��F<��<#3�<s�<�{�<��<#3�<��<��F<��;��U�NzV���%�
��X.�
kF�H�N�.kF��X.��
���pzV���U�`   `   1��;@�_<6Y�<�U�<��<��<�U�<WY�<s�_<��;��Q��+�ف�����X.���N��$`�|$`��N�Y.���́���+���Q�`   `   ' <[�z<�M�<k8�<��<k8�<�M�<\�z< <pr ;��׻%����R�` �
kF��$`�EAi��$`�kF�` ��R�%�����׻or ;`   `   �J<y1�<��<\��<���<��<S1�<zJ<���;���x;������F}/�H�N�|$`��$`�W�N�5}/�������x;����9��;`   `   ��q<m�<d�<
h�<�<m�<�q<�i<"�B;ʫ�וp��ʼ���5}/�-kF��N�kF�5}/�Ё��ʼ��p�ʫ���B;�i<`   `   ��<�d�<[Q�<{Q�<�d�<��<YQT<Q�;��o:~��;���<�ʼ��` ��X.�Y.�` ����ʼ4���ף�n�o:Q�;�QT<`   `   �ח<�<�Y�<�<�ח<�!�<L�@<G2�;�`F9ף�f�p����S����
����R������p�ף滒xF9G2�;��@<�!�<`   `   �k�<���<j��<�k�<�v�<Ȱx<N�9<�2�;��o:�ʫ��x;�����ف��+����́��$����x;�ʫ�q�o:G2�;��9<ϰx<�v�<`   `   ���<혬<(��<���<��<ϰx<�@<Q�;�B;���V�׻�+�zV�<xe�ozV��+���׻�����B;Q�;��@<ϰx<�<���<`   `   )��<��<���<���<�v�<�!�<YQT<�i<���;�s ;��Q�w�U�s���>�����U���Q�qr ;9��;�i<�QT<�!�<�v�<���<���<`   `   [X�<Z��<���<���<_ʹ<�8�<2�<�<H�<��<k\�<H��<"�<H��<T\�<��<n�<�<�1�<�8�<�ʹ<���<p��<Z��<`   `   Z��<�V�<x��<U3�<�(�<�(�<�<�+�<�٧<�ע< �<i̜<f̜<	�<�ע<z٧<�+�<#�<�(�<�(�<L3�<���<V�<K��<`   `   ���<x��<�N�<��<�E�<C˽<r�<|X�<�ط<lu�<�<��<�<lu�<�ط<|X�<r�<C˽<�E�<��<�N�<x��<���<�Ļ<`   `   ���<T3�<��<d��<�u�<�I�<�=�<�^�<���<J�<���<��<J�<���<�^�<�=�<uI�<nu�<t��<��<L3�<���<�ͷ<�ͷ<`   `   _ʹ<�(�<�E�<�u�<�(�<���<`��<���<�{�<���<x��<���<�{�<���<7��<���<)�<�u�<�E�<�(�<wʹ<aر<�ϰ<aر<`   `   �8�<�(�<C˽<�I�<���<���<���<V��<�S�<+�<+�<�S�<R��<į�<���<���<tI�<\˽<�(�<�8�<��<���<���<��<`   `   2�<�<r�<�=�<`��<���<k��<�y�<��<rH�<���<�y�<R��<���<q��<�=�<r�<�<2�<6�<�V�<�g�<�V�<6�<`   `   �<�+�<|X�<�^�<���<V��<�y�<>b�<wS�<bS�<5b�<�y�<R��<f��<�^�<�X�<�+�<
�<�<�$�<�Q�<�Q�<�$�<�<`   `   G�<�٧<�ط<���<�{�<�S�<��<wS�<��<wS�<l��<�S�<�{�<���<�ط<�٧<i�<�0�<7t<9�b<Fy\<8�b<]t<�0�<`   `   ��<�ע<ku�<J�<���<+�<rH�<bS�<wS�<�H�<+�<��<J�<�u�<�ע<	��<�t<)@P<$�4<0&<&<�4<$@P<�t<`   `   j\�<��<�<���<x��<+�<���<5b�<l��<+�<���<���<ݷ�< �<l\�<HG]<QF.<V*<�H�;���;�H�;V*<2F.<HG]<`   `   H��<i̜<��<��<���<�S�<�y�<�y�<�S�<��<���<�<e̜<9��<j�K<I<�g�;jB[;��;X�;#B[;Bh�;D<O�K<`   `   !�<e̜<�<J�<�{�<R��<R��<R��<�{�<J�<ݷ�<e̜<4�<c=B<�~�;^�|;��:z~Ӻ9�z~Ӻ��:^�|;�~�;c=B<`   `   H��<	�<ku�<���<���<į�<���<f��<���<�u�< �<9��<c=B<CJ�;�<9;h����;��Y�ǻ�ǻm;������-<9;8J�;j=B<`   `   T\�<�ע<�ط<�^�<7��<���<q��<�^�<�ط<�ע<l\�<j�K<�~�;�<9;����y���w���3����z���$����<9;�~�;j�K<`   `   ��<z٧<|X�<�=�<���<���<�=�<�X�<�٧<	��<IG]<J<`�|;f���y���V�i�:�E�:�5���������z�|;D<[G]<`   `   n�<�+�<r�<tI�<)�<tI�<r�<�+�<i�<�t<QF.<�g�;��:�;��w��i�:�gK�i�:�}���;��}�:�g�;DF.<�t<`   `   �<#�<C˽<nu�<�u�<\˽<�<
�<�0�<*@P<W*<mB[;t~ӺX�ǻ�3�D�:�i�:��3��ǻ@~Ӻ&B[;i*<$@P<�0�<`   `   �1�<�(�<�E�<t��<�E�<�(�<2�<�<8t<%�4<�H�;��;9��ǻ���5�}���ǻ�9���;�H�;%�4<ft<�<`   `   �8�<�(�<��<��<�(�<�8�<6�<�$�<9�b<1&<���;\�;r~Ӻk;��x��������;��>~Ӻ��;��;&<�b<�$�<R�<`   `   �ʹ<L3�<�N�<L3�<wʹ<��<�V�<�Q�<Gy\<&<�H�;'B[;��:𾦺���𾦺��:'B[;�H�;&<�y\<�Q�<rV�<��<`   `   ���<���<x��<���<aر<���<�g�<�Q�<9�b<�4<W*<Dh�;b�|;1<9;�<9;|�|;�g�;i*<%�4<�b<�Q�<�g�<���<Cر<`   `   p��<V�<���<�ͷ<�ϰ<���<�V�<�$�<^t<%@P<3F.<E<�~�;9J�;�~�;E<EF.<%@P<gt<�$�<sV�<���<�ϰ<�ͷ<`   `   Z��<K��<�Ļ<�ͷ<aر<��<6�<�<�0�<�t<IG]<P�K<d=B<k=B<k�K<[G]<�t<�0�<�<R�<��<Cر<�ͷ<�Ļ<`   `   �<3��<��<�/�<�w�<�i�<���<���<X��<�}�<��<�3�<���<�3�<��<�}�<g��<���<���<�i�<�w�<�/�<ܨ�<3��<`   `   3��<�,�<��<Z��<^�<��<�E�<���<���<���<���<���<���<���<���<���<���<�E�<��<^�<]��<(��<�,�<'��<`   `   ��<��<���<�Y�<��<v�<���<�]�<Jt�<�U�<�1�<p �<�1�<�U�<Zt�<�]�<���<v�<.��<�Y�<���<��<���<^Z�<`   `   �/�<Z��<�Y�<���<�m�<ٞ�<�W�<u��<�E�<���<��<��<���<rE�<t��<�W�<؞�<�m�<���<�Y�<]��<�/�<�,�<�,�<`   `   �w�<^�<��<�m�<|��<���<�&�<���<���<�w�<��<�w�<���<���<~&�<���<���<�m�<��<^�<�w�<��<��<��<`   `   �i�<��<v�<ٞ�<���<zX�<|�<��<�H�<���<���<�H�<��<��<yX�<���<؞�<��<��<�i�<N�<ٜ�<ќ�<N�<`   `   ���<�E�<���<�W�<�&�<|�<�"�<�3�<I`�<o��<b`�<�3�<�"�<|�<�&�<�W�<���<�E�<���<�~�<y��<k��<���<�~�<`   `   ���<���<�]�<u��<���<��<�3�<G<�<1A�<"A�<=<�<4�<��<r��<t��<�]�<���<���<��<Ρ�<�>�<�>�<ơ�<��<`   `   X��<���<Jt�<�E�<���<�H�<I`�<1A�<:��<1A�<B`�<�H�<���<�E�<;t�<���<e��<I4�<��<<׮<�g�<<׮<"��<I4�<`   `   �}�<���<�U�<���<�w�<���<o��<"A�<1A�<���<���<�w�<���<�U�<���<�}�<7�<��<D��<�\�<�\�<D��<��<7�<`   `   ��<���<�1�<��<��<���<b`�<=<�<B`�<���<���<��<�1�<���<��<���<.�<8��<�ʘ<QƖ<�ʘ<8��<.�<���<`   `   �3�<���<p �<��<�w�<�H�<�3�<4�<�H�<�w�<��<� �<���<~3�<9ͮ<X�<	+�<d��<��<��<g��<	+�<�W�<:ͮ<`   `   ���<���<�1�<���<���<��<�"�<��<���<���<�1�<���<��<�H�<`�<㎑<;=�<^`}<�x<^`}<7=�<⎑<g�<�H�<`   `   �3�<���<�U�<qE�<���<��<|�<r��<�E�<�U�<���<~3�<�H�<���<M��<~��<U�k<�}`<�}`<W�k<���<N��<y��<{H�<`   `   ��<���<Yt�<t��<}&�<yX�<�&�<t��<;t�<���<��<9ͮ<`�<M��<;<}<��b<*�P<�vJ<)�P<��b<3<}<M��<m�<9ͮ<`   `   �}�<���<�]�<�W�<���<���<�W�<�]�<���<�}�<���<X�<㎑<~��<��b<�/K<��><��><�/K<��b<���<ގ�<�W�<���<`   `   g��<���<���<؞�<���<؞�<���<���<e��<7�<.�<	+�<;=�<V�k<+�P<��><68<��><(�P<V�k<==�<	+�<.�<7�<`   `   ���<�E�<v�<�m�<�m�<��<�E�<���<I4�<��<9��<d��<_`}<�}`<�vJ<��><��><�vJ<�}`<U`}<g��<B��<��<:4�<`   `   ���<��<.��<���<��<��<���<��<��<D��<�ʘ<��<�x<�}`<)�P<�/K<)�P<�}`<�x<��<{ʘ<D��<1��<��<`   `   �i�<^�<�Y�<�Y�<^�<�i�<�~�<Ρ�<=׮<�\�<RƖ<��<_`}<W�k<��b<��b<V�k<U`}<��<\Ɩ<�\�<.׮<ǡ�<�~�<`   `   �w�<]��<���<]��<�w�<N�<z��<�>�<�g�<�\�<�ʘ<g��<8=�<���<3<}<���<==�<g��<{ʘ<�\�<�g�<�>�<p��<N�<`   `   �/�<(��<��<�/�<��<ٜ�<k��<�>�<=׮<E��<9��<
+�<㎑<N��<M��<ގ�<	+�<C��<E��<.׮<�>�<}��<ќ�<���<`   `   ܨ�<�,�<���<�,�<��<ќ�<���<ǡ�<#��<��<.�<�W�<g�<y��<m�<�W�<.�<��<1��<ǡ�<p��<ќ�<3��<�,�<`   `   3��<'��<^Z�<�,�<��<N�<�~�<��<I4�<7�<���<:ͮ<�H�<{H�<9ͮ<���<7�<;4�<��<�~�<N�<���<�,�<oZ�<`   `   ���<A'�<ǣ�<hb�<zY�<�q�<�<���<��<�f�<��<�B�<�]�<�B�<��<�f�<��<���<˖�<�q�<sY�<hb�<ˣ�<A'�<`   `   A'�<X��<%��<z��<A�<���<�O�<&��<\��<O��<Ԁ�<'��<2��<݀�<B��<U��<4��<�O�<���<A�<���<+��<M��<9'�<`   `   ǣ�<%��<r��<Ӳ�<��<�z�<�@�<���<��<s	�<���<���<s��<s	�<�<���<�@�<�z�<*��<Ӳ�<_��<%��<ڣ�<�K�<`   `   hb�<z��<Ӳ�<G��<��< >�<�&�<ƻ�<���<���<$1�<-1�<���<���<���<�&�<>�<��<9��<ڲ�<���<`b�<��<��<`   `   zY�<A�<��<��<v��<���<���<�H�<_Y�<���<5�<���<[Y�<�H�<���<���<m��<��<��<A�<vY�<��<��<��<`   `   �q�<���<�z�< >�<���<�#�<%��<�Y�<9�<���<���<9�<�Y�<*��<�#�<���<>�<�z�<���<�q�<���<&��<��<���<`   `   �<�O�<�@�<�&�<���<%��<*��<N��<r��<���<���<N��<��<%��<���<�&�<�@�<�O�<ٖ�<�h�<���<�y�<��<�h�<`   `   ���<%��<���<ƻ�<�H�<�Y�<N��<���<|J�<uJ�<���<S��<�Y�<�H�<���<���<3��<~��<a�<��<�	�<�	�<��<n�<`   `   ��<\��<��<���<_Y�<9�<r��<|J�<���<|J�<u��<9�<YY�<���<��<\��<��<���<?�<[e�<���<[e�<<�<���<`   `   �f�<O��<s	�<���<���<���<���<uJ�<|J�<���<���<���<���<y	�<B��<�f�<���<���<���<E�<!E�<���<���<���<`   `   ��<Ԁ�<���<$1�<5�<���<���<���<u��<���<!5�<$1�<u��<Ԁ�<+��<�+�<���<���<�z�<���<�z�<���<���<�+�<`   `   �B�<'��<���<-1�<���<9�<N��<S��<9�<���<$1�<���<2��<�B�<�D�<�0�<�z�<d��<y�<��<p��<�z�<�0�<�D�<`   `   �]�<2��<r��<���<[Y�<�Y�<��<�Y�<YY�<���<u��<2��<�]�<�M�<L��<`��<~�<��<Գ�<��<��<`��<J��<�M�<`   `   �B�<݀�<s	�<���<�H�<*��<%��<�H�<���<y	�<Ԁ�<�B�<�M�<9��<j(�<w��<9��<$��<��<+��<���<w(�<.��<�M�<`   `   ��<B��<�<���<���<�#�<���<���<��<B��<+��<�D�<L��<j(�<�z�<K}�<���<nֿ<���<K}�<iz�<j(�<b��<�D�<`   `   �f�<U��<���<�&�<���<���<�&�<���<\��<�f�<�+�<�0�<`��<w��<K}�<}�<�8�<�8�<o�<X}�<���<U��<�0�<�+�<`   `   ��<3��<�@�<>�<m��<>�<�@�<3��<��<���<���<�z�<~�<9��<���<�8�<tQ�<�8�<���<9��<}�<�z�<���<���<`   `   ���<�O�<�z�<��<��<�z�<�O�<~��<���<���<���<d��<��<$��<nֿ<�8�<�8�<{ֿ<��<t��<p��<���<���<���<`   `   ˖�<���<*��<9��<��<���<ٖ�<a�<?�<���<�z�<y�<Գ�<��<���<o�<���<��<��<y�<�z�<���<Q�<a�<`   `   �q�<A�<Ӳ�<ڲ�<A�<�q�<�h�<��<\e�<E�<���<��<��<+��<L}�<Y}�<9��<t��<y�<��<!E�<Ue�<��<�h�<`   `   sY�<���<_��<���<vY�<���<���<�	�<���<!E�<�z�<p��<��<���<iz�<���<}�<p��<�z�<!E�<���<�	�<���<���<`   `   hb�<+��<%��<`b�<��<&��<�y�<�	�<\e�<���<���<�z�<`��<w(�<j(�<U��<�z�<���<���<Ue�<�	�<�y�<��<��<`   `   ˣ�<M��<ڣ�<��<���<��<��<��<<�<���<���<�0�<J��</��<b��<�0�<���<���<Q�<��<���<��<���<��<`   `   A'�<9'�<�K�<��<��<���<�h�<o�<���<���<�+�<�D�<�M�<�M�<�D�<�+�<���<���<a�<�h�<���<��<��<�K�<`   `   ��<d�<�%�<k\�<X��<���<��<�@�<�a�< D�<���<���<z�<���<���< D�<�a�<�@�<��<���<=��<k\�<�%�<d�<`   `   d�<���<s��<
f�<.�<1�<�T�<Hj�<V�<���<��<8��<G��<��<���<V�<aj�<�T�<�0�<.�<f�<p��<���<d�<`   `   �%�<s��<�6�<z��<��<��<���<���<ZI�<��<a�<*��<�`�<��<oI�<���<��<��<-��<z��<6�<s��<�%�<���<`   `   k\�<
f�<z��<H��<+x�<�a�<]3�<���<�(�<#�<���<���<2�<�(�<���<V3�<�a�<3x�</��<v��<f�<h\�<���<��<`   `   X��<.�<��<+x�<�D�<��<���<7��<
��<���<9��<���<���<7��<���<��<�D�<+x�<8��<.�<G��<!9�<2��<!9�<`   `   ���<1�<��<�a�<��<��<���<��<s�<P��<J��<s�<��<���<��<��<�a�<��<�0�<���<���<#�<�<���<`   `   ��<�T�<���<]3�<���<���<ڹ�<�l�<K��<Q�<P��<�l�<ѹ�<���<���<]3�<��<�T�<��</�<|a�<�(�<�a�</�<`   `   �@�<Gj�<���<���<7��<��<�l�<}��<�<�<w��<�l�<��<>��<���<���<aj�<�@�</A�<���< $�<$�<���<HA�<`   `   �a�<V�<ZI�<�(�<
��<s�<K��<�<T�<�<X��<s�<���<�(�<tI�<V�<�a�<��<���<�N�<$�<�N�<���<��<`   `    D�<���<��<#�<���<P��<Q�<�<�<K�<J��<���<2�< ��<���<�C�<I��<d��<y�<�4�<�4�<5y�<X��</��<`   `   ���<��<a�<���<9��<J��<P��<w��<X��<J��<8��<���<�`�<��<���<9Q�<���<�s�<�)�<��<�)�<�s�<���<9Q�<`   `   ���<8��<*��<���<���<s�<�l�<�l�<s�<���<���<&��<G��<}��<;��<�Y�<��<���<Ұ�<��<���<��<�Y�<Q��<`   `   z�<G��<�`�<2�<���<��<ѹ�<��<���<2�<�`�<G��<n�<A7�<
K�<>�<��<Q��<O��<P��<��<>�< K�<A7�<`   `   ���<��<��<�(�<7��<���<���<>��<�(�< ��<��<}��<A7�<��<���<l��<���<��<���<���<���<���<���<27�<`   `   ���<���<oI�<���<���<��<���<���<tI�<���<���<;��<
K�<���<+�<T�<�`�<�b�<�`�<T�<�*�<���<%K�<;��<`   `    D�<V�<���<V3�<��<��<]3�<���<V�<�C�<9Q�<�Y�<>�<l��<T�<��<���<s��<���<,T�<���<>�<�Y�<?Q�<`   `   �a�<aj�<��<�a�<�D�<�a�<��<aj�<�a�<I��<���<��<��<���<�`�<���<��<���<�`�<���<��<��<���<I��<`   `   �@�<�T�<��<2x�<+x�<��<�T�<�@�<��<d��<�s�<���<Q��<��<�b�<s��<���<�b�<���<A��<���<�s�<X��<��<`   `   ��<�0�<-��</��<8��<�0�<��</A�<���<y�<�)�<Ұ�<O��<���<�`�<���<�`�<���<x��<Ұ�<�)�<y�<���</A�<`   `   ���<.�<z��<v��<.�<���</�<���<�N�<�4�<��<��<Q��<���<T�<,T�<���<A��<Ұ�<��<�4�<�N�<���<)�<`   `   =��<f�<6�<f�<H��<���<|a�< $�<$�<�4�<�)�<���<��<���<�*�<���<��<���<�)�<�4�<�#�< $�<�a�<���<`   `   k\�<p��<s��<h\�<!9�<#�<�(�<$�<�N�<5y�<�s�<��<>�<���<���<>�<��<�s�<y�<�N�< $�<�(�<�<(9�<`   `   �%�<���<�%�<���<2��<�<�a�<���<���<Y��<���<�Y�< K�<���<%K�<�Y�<���<Y��<���<���<�a�<�<6��<���<`   `   d�<d�<���<��<!9�<���</�<HA�<��</��<9Q�<Q��<A7�<27�<;��<@Q�<I��<��</A�<)�<���<(9�<���<���<`   `   ��<R�<��<�N�<B��<��<�K�<��<:��<��<2��<���<��<���<K��<��<��<��</L�<��<��<�N�<��<R�<`   `   R�<P��<t��<��<I��<���<U��<��<\��<w��<���<;j�<Lj�<���<Z��<f��<5��<C��<���<\��<�<f��<E��<R�<`   `   ��<t��<��<�<���<���<�}�<rK�<��<�#�<{��<6�<g��<�#�<��<rK�<�}�<���<��<�<߶�<t��<��<��<`   `   �N�<��<�<�p�<���<��<�,�<��<���<��<�.�<�.�< ��<���<š�<�,�<;��< ��<rp�<�<�<�N�<���<���<`   `   B��<H��<���<���<�C�<I��<H��<���<���<A_�<s��<A_�<}��<���<v��<I��<�C�<���<%��<H��<'��<m��<�V�<m��<`   `   ��<���<���<��<I��<���<d~�<-E�<���<��<��<���<>E�<R~�<���<]��<;��<���<���<��<��<�B�<�B�<˃�<`   `   �K�<T��<�}�<�,�<H��<d~�<6�<F��<���<���<���<F��<7�<d~�<Q��<�,�<�}�<T��<L�<���<���<g��<Ӝ�<���<`   `   ��<��<rK�<��<���<-E�<F��<��<z��<���<��<4��<>E�<���<š�<dK�<4��<��<�r�<�H�<�1�<�1�<�H�<�r�<`   `   :��<\��<��<���<���<���<���<z��<s��<z��<��<���<s��<���<-��<\��<��<S�<,�<Z�<�"�<Z�<�<S�<`   `   ��<w��<�#�<��<A_�<��<���<���<z��<���<��<T_�< ��<�#�<Z��<��<�{�<��<z�<�>�<�>�<��<���<�{�<`   `   1��<���<{��<�.�<s��<��<���<��<��<��<c��<�.�<w��<���<K��<Ȋ�<.P�<���<�N�<�p�<IN�<���<\P�<Ȋ�<`   `   ���<;j�<6�<�.�<A_�<���<F��<4��<���<T_�<�.�<6�<Lj�<���<�	�<3E�<�M�<�<�m�<�m�<��<�M�<'E�<
�<`   `   ��<Lj�<f��< ��<}��<>E�<7�<>E�<s��< ��<w��<Lj�<��<V��<=��<r�<�3�<p��<�0�<p��<�3�<r�<,��<V��<`   `   ���<���<�#�<���<���<R~�<d~�<���<���<�#�<���<���<V��<���<��<V��<���<�\�<�\�<���<o��<2��<���<E��<`   `   K��<Z��<��<š�<v��<���<Q��<š�<-��<Z��<L��<�	�<=��<��<@�<R��<#��<��<e��<R��<�<��<Y��<�	�<`   `   ��<e��<rK�<�,�<I��<]��<�,�<dK�<\��<��<Ȋ�<3E�<r�<V��<R��<�9�<N�<,�<�9�<n��<o��<a�<'E�<ˊ�<`   `   ��<4��<�}�<;��<�C�<;��<�}�<4��<��<�{�<.P�<�M�<�3�<���<#��<N�<�u�<N�<'��<���<�3�<�M�<7P�<�{�<`   `   ��<C��<���< ��<���<���<U��<��<S�<��<���<�<p��<�\�<��<,�<N�<��<�\�<_��<��<���<���<]�<`   `   /L�<���<��<rp�<%��<���<L�<�r�<,�<z�<�N�<�m�<�0�<�\�<e��<�9�<'��<�\�<�0�<�m�<gN�<z�<.�<�r�<`   `   ��<\��<�<�<I��<��<���<�H�<Z�<�>�<�p�<�m�<p��<���<R��<n��<���<_��<�m�<�p�<�>�<c�<�H�<r��<`   `   ��<�<߶�<�<'��<��<���<�1�<�"�<�>�<IN�<��<�3�<o��<�<o��<�3�<��<gN�<�>�<�"�<�1�<͜�<��<`   `   �N�<f��<t��<�N�<m��<�B�<g��<�1�<Z�<��<���<�M�<r�<3��<��<a�<�M�<���<z�<c�<�1�<U��<�B�<���<`   `   ��<E��<��<���<�V�<�B�<Ԝ�<�H�<�<���<\P�<'E�<,��<���<Y��<'E�<7P�<���<.�<�H�<͜�<�B�<�V�<���<`   `   R�<R�<��<���<m��<˃�<���<�r�<S�<�{�<Ȋ�<
�<V��<E��<�	�<ˊ�<�{�<]�<�r�<r��<��<���<���<��<`   `   .�<d=�<*��<��<�a�<�-�<|4�<�V�<�i�<TB�<���<���<���<���<ݷ�<TB�<di�<�V�<�4�<�-�<Va�<��<K��<d=�<`   `   d=�<ӟ�<�`�<�x�<:��<���<!l�<�D�<[��<�p�<h}�<x
�<�
�<g}�<�p�<m��<E�<l�<v��<X��<�x�<�`�<ʟ�<l=�<`   `   *��<�`�<�2�<�G�<9��< �<���<�9�<t��<��<FU�<&��<6U�<��<���<�9�<���< �<@��<�G�<�2�<�`�<,��<��<`   `   ��<�x�<�G�<~Q�<�y�<���<��<�8�<(9�<��<nS�<mS�<'��<:9�<�8�<e�<Ͽ�<�y�<YQ�<�G�<�x�<��<Z��<d��<`   `   �a�<:��<9��<�y�<2i�<�n�<�e�<�B�<f��<E`�<���<E`�<D��<�B�<�e�<�n�<�h�<�y�<u��<:��<la�<��<���<��<`   `   �-�<���< �<���<�n�<
&�<x��<�U�<���<���<���<���<�U�<[��<�%�<�n�<Ͽ�<��<v��<�-�<A��<��<	��<&��<`   `   |4�<!l�<���<��<�e�<x��<�(�<Yt�<:��<��<'��<Yt�<�(�<x��<�e�<��<}��<!l�<�4�<{�<���<���<���<{�<`   `   �V�<�D�<�9�<�8�<�B�<�U�<Yt�<���<��<��<���<=t�<�U�<�B�<�8�<�9�<E�<�V�<ri�<�y�<,��<��<�y�<�i�<`   `   �i�<[��<t��<(9�<f��<���<:��<��<��<��<U��<���<7��<(9�<���<[��<mi�<���<n�<�S�<.f�<�S�<S�<���<`   `   TB�<�p�<��<��<E`�<���<��<��<��<��<���<c`�<'��<���<�p�<\B�<�	�<��<,1�<=s�<Ws�<Q1�<���<m	�<`   `   ���<h}�<FU�<nS�<���<���<'��<���<U��<���<���<nS�<LU�<h}�<ӷ�<}��<8�<���<�p�<���<�p�<���<h�<}��<`   `   ���<x
�<&��<mS�<E`�<���<Yt�<=t�<���<c`�<nS�<��<�
�<§�<M�<��<*�<��<E��<j��<��<�)�<��<5M�<`   `   ���<�
�<6U�<'��<D��<�U�<�(�<�U�<7��<'��<LU�<�
�<���<B�<��<'��<4<�<�#�<�r�<�#�<A<�<'��<��<B�<`   `   ���<g}�<��<:9�<�B�<[��<x��<�B�<(9�<���<h}�<§�<B�<�o�<(��<t��<���<���<���<���<���<H��<�o�<1�<`   `   ܷ�<�p�<���<�8�<�e�<�%�<�e�<�8�<���<�p�<ӷ�<M�<��<(��<7�<���<�%�<ϑ�<I&�<���<��<(��<��<M�<`   `   TB�<m��<�9�<e�<�n�<�n�<��<�9�<[��<\B�<}��<��<'��<t��<���<��<܎�<���<ݦ�<��<���<��<��<|��<`   `   di�<E�<���<Ͽ�<�h�<Ͽ�<}��<E�<mi�<�	�<8�<*�<5<�<���<�%�<܎�<��<܎�<&�<���<+<�<*�<C�<�	�<`   `   �V�<l�< �<�y�<�y�<��<!l�<�V�<���<��<���<��<�#�<���<ϑ�<���<܎�<��<���<�#�<��<���<���<���<`   `   �4�<v��<@��<YQ�<u��<v��<�4�<ri�<n�<,1�<�p�<E��<�r�<���<I&�<ݦ�<&�<���<s�<E��<�p�<,1�<g�<ri�<`   `   �-�<X��<�G�<�G�<:��<�-�<{�<�y�<�S�<=s�<���<j��<�#�<���<���<��<���<�#�<E��<���<Ws�<�S�<�y�<_�<`   `   Va�<�x�<�2�<�x�<ma�<A��<���<,��<.f�<Ws�<�p�<��<A<�<���<��<���<+<�<��<�p�<Ws�<f�<,��<���<A��<`   `   ��<�`�<�`�<��<��<��<���<��<�S�<Q1�<���<�)�<'��<H��<(��<��<*�<���<,1�<�S�<,��<g��<
��<�<`   `   K��<ʟ�<,��<Z��<���<
��<���<�y�<S�<���<h�<��<��<�o�<��<��<C�<���<g�<�y�<���<
��<���<Z��<`   `   d=�<l=�<��<d��<��<&��<{�<�i�<���<m	�<}��<6M�<B�<1�<M�<|��<�	�<���<ri�<_�<A��<�<Z��<��<`   `   ;�<�K�<���<ٮ�<���<}G�<���</��<�P�<���<���<��<��<��< �<���<ZP�</��<��<}G�<A��<ٮ�<���<�K�<`   `   �K�<���<�5�<��<�=�<���<��<*y�<���<`�<���<�I�<	J�<���<@�<���<Ry�<n�<ԍ�<
>�<��<�5�<���<
L�<`   `   ���<�5�<2��<@��<���<X��<a$�<�U�<he�<�<�<��<���<��<�<�<oe�<�U�<]$�<X��<���<@��<6��<�5�<���<��<`   `   ٮ�<��<@��<�|�<�d�<n\�<�R�<�<�<d�<ؐ�<C��<>��<��<}�<�<�<�R�<�\�<�d�<�|�<"��<��<��<�w�<�w�<`   `   ���<�=�<���<�d�<P�<���<���<'5�<��<��<4#�<��<Ƶ�<'5�<:��<���< �<�d�<��<�=�<Z��<���<f��<���<`   `   }G�<���<X��<n\�<���<U�<���<�3�<��<��<��<��<�3�<���<�T�<���<�\�<9��<ԍ�<�G�<��<�<�<��<`   `   ���<��<a$�<�R�<���<���<��<�9�<8[�<�f�<[�<�9�<��<���<��<�R�<V$�<��<���<���<���<���<���<���<`   `   /��<)y�<�U�<�<�<'5�<�3�<�9�<�A�<G�<!G�<�A�<�9�<�3�<N5�<�<�<bU�<Ry�<=��<r��<z��<��<���<s��<���<`   `   �P�<���<he�<d�<��<��<8[�<G�<�?�<G�<W[�<��<���<d�<�e�<���<eP�<���<��<�W�<�l�<�W�<��<���<`   `   ���<`�<�<�<א�<��<��<�f�<!G�<G�<yf�<��<�<��<w<�<@�<���<���<�@�<���<N �<h �<��<�@�<͕�<`   `   ���<���<��<C��<4#�<��<[�<�A�<W[�<��<#�<C��<,��<���< �<1$�<�+�<���<7��<���<���<���<�+�<1$�<`   `   ��<�I�<���<>��<��<��<�9�<�9�<��<�<C��<���<J�<��<DD�<��<6��<���<g;�<�;�<���<��<��<dD�<`   `   ��<J�<��<��<Ƶ�<�3�<��<�3�<���<��<,��<J�<��<���<���<�E�<���<6^�<g��<6^�<���<�E�<��<���<`   `   ��<���<�<�<}�<'5�<���<���<N5�<d�<w<�<���<��<���<���<��<\��<q��<���<y��<H��<v��<4��<���<|��<`   `    �<@�<oe�<�<�<:��<�T�<��<�<�<�e�<@�< �<DD�<���<��<,�<��<��<�+�<i��<��<��<��<��<DD�<`   `   ���<���<�U�<�R�<���<���<�R�<bU�<���<���<1$�<��<�E�<\��<��<�:�<��<g�<�:�<4��<v��<�E�<��<,$�<`   `   ZP�<Ry�<]$�<�\�< �<�\�<V$�<Ry�<eP�<���<�+�<6��<���<q��<��<��<Yo�<��< ��<q��<���<6��<�+�<���<`   `   /��<n�<X��<�d�<�d�<9��<��<=��<���<�@�<���<���<6^�<���<�+�<g�<��<�+�<y��<'^�<���<���<�@�<���<`   `   ��<ԍ�<���<�|�<��<ԍ�<���<r��<��<���<7��<g;�<h��<y��<i��<�:�< ��<y��<���<g;�<"��<���<��<r��<`   `   }G�<
>�<@��<"��<�=�<�G�<���<z��<�W�<N �<���<�;�<6^�<H��<��<4��<q��<'^�<g;�<���<h �<X�<s��<���<`   `   A��<��<6��<��<Z��<��<���<��<�l�<h �<���<���<���<v��<��<v��<���<���<"��<h �<�l�<��<���<��<`   `   ٮ�<�5�<�5�<��<���<�<���<���<�W�<��<���<��<�E�<4��<��<�E�<6��<���<���<X�<��<u��<�<���<`   `   ���<���<���<�w�<f��<�<���<s��<��<�@�<�+�<��<��<���<��<��<�+�<�@�<��<s��<���<�<F��<�w�<`   `   �K�<
L�<��<�w�<���<��<���<���<���<͕�<1$�<dD�<���<|��<DD�<,$�<���<���<r��<���<��<���<�w�<��<`   `   ���<���<��<���<���<��<��<�]�<y��<���<U��<nF�<�y�<nF�<}��<���<3��<�]�<�<��<K��<���<��<���<`   `   ���<��<�b�<��<���<� �<��<�;�<3B�<#�<���<L�<Y�<���<�"�<QB�<<�<��<� �<"��<��<�b�<{��<���<`   `   ��<�b�<m��<��<�[�<SA�<�1�<��<>��<���<���<�<���<���<@��<��<�1�<SA�<�[�<��<x��<�b�<��<���<`   `   ���<��<��<�$�<��<���<�L�<W��<B��<!��<�2�<�2�<.��<_��<8��<�L�<��<I��<�$�<Ό�<��<���<֙�<ڙ�<`   `   ���<���<�[�<��<Y�<$��<o�<4��<tI�<���<̜�<���<JI�<4��<[o�<$��<�X�<��<�[�<���<f��<���<�t�<���<`   `   ��<� �<SA�<���<$��<�@�<v��<9��<��<�1�<�1�<��<E��<K��<x@�<Q��<��</A�<� �<��<���<���<���<���<`   `   ��<��<�1�<�L�<o�<v��<���<t��< ��<��<���<t��<���<v��<o�<�L�<�1�<��<��<C�<��<�<�<C�<`   `   �]�<�;�<��<V��<4��<9��<t��<S��<b��<���<]��<J��<E��<a��<8��<��<<�<�]�<e��<���<��< ��<���<���<`   `   y��<3B�<>��<A��<tI�<��< ��<b��<	��<b��<A��<��<:I�<A��<���<3B�<?��<i�<UP�<��<���<��<4P�<i�<`   `   ���<#�<���<!��<���<�1�<��<���<b��<���<�1�<҇�<.��<b��<�"�<���<�l�<d��<�]�<���<ѓ�<^�<`��<hl�<`   `   U��<���<���<�2�<̜�<�1�<���<]��<A��<�1�<���<�2�<���<���<b��<���<Lq�<��<n��<��<0��<��<xq�<���<`   `   nF�<L�<�<�2�<���<��<t��<J��<��<҇�<�2�<��<Y�<�F�<[y�<w��<��<�F�< ��<&��<G�<ʒ�<s��<yy�<`   `   �y�<Y�<���<.��<JI�<E��<���<E��<:I�<.��<���<Y�<ry�<Z��<�Z�<g��<ը�<�O�<Q��<�O�<��<g��<�Z�<Z��<`   `   nF�<���<���<_��<4��<K��<v��<a��<A��<b��<���<�F�<Z��<Q��<X3�<���<���<	�<��<���<��<w3�<M��<M��<`   `   }��<�"�<@��<8��<[o�<x@�<o�<8��<���<�"�<b��<[y�<�Z�<X3�<���<�'�<���<�H�<9��<�'�<h��<X3�<�Z�<[y�<`   `   ���<QB�<��<�L�<$��<Q��<�L�<��<3B�<���<���<w��<g��<���<�'�<,S�<���<i��<S�<�'�<��<Z��<s��<w��<`   `   3��<<�<�1�<��<�X�<��<�1�<<�<?��<�l�<Lq�<��<ը�<���<���<���<BE�<���<���<���<ʨ�<��<Yq�<�l�<`   `   �]�<��<SA�<I��<��</A�<��<�]�<i�<d��<��<�F�<�O�<	�<�H�<i��<���<�H�<��<�O�<G�<��<`��<��<`   `   �<� �<�[�<�$�<�[�<� �<��<e��<UP�<�]�<n��<��<Q��<��<9��<S�<���<��<���<��<_��<�]�<<P�<e��<`   `   ��<"��<��<Ό�<���<��<C�<���<��<���<��<&��<�O�<���<�'�<�'�<���<�O�<��<��<ѓ�<.��<���<�<`   `   K��<��<x��<��<f��<���<��<��<���<ғ�<0��<G�<��<��<h��<��<ʨ�<G�<_��<ѓ�<b��<��<�<���<`   `   ���<�b�<�b�<���<���<���<�< ��<��<^�<��<ʒ�<g��<w3�<X3�<Z��<��<��<�]�<.��<��<��<���<�<`   `   ��<{��<��<֙�<�t�<���<�<���<4P�<`��<xq�<s��<�Z�<M��<�Z�<s��<Yq�<`��<<P�<���<�<���<�t�<֙�<`   `   ���<���<���<ڙ�<���<���<C�<���<i�<hl�<���<yy�<Z��<N��<[y�<w��<�l�<��<e��<�<���<�<֙�<���<`   `   n\�<Ly�<���<�V�<��<���<��<���<d��<���<�Y�<:��<���<:��<Z�<���<��<���<S��<���<K�<�V�<��<Ly�<`   `   Ly�<%��<W
�<��<�D�<��<���<��<<��<�.�<���<��<!��<��<�.�<\��<��<i��<h�<�D�<#��<1
�<$��<ay�<`   `   ���<W
�<�l�<��<���<�<�<���<���<�9�<���<- �<��</ �<���<�9�<���<���<�<�<���<��<�l�<W
�<���<]��<`   `   �V�<��<��<c�<���<�t�<�<���<F��<C�<2m�<&m�< C�<g��<���<��<�t�<���<�b�<���<#��<�V�<�6�<�6�<`   `   ��<�D�<���<���<&K�<e��<��<�r�<߸�<���<���<���<���<�r�<�<e��<�J�<���<��<�D�<f�<Z��<���<Z��<`   `   ���<��<�<�<�t�<e��<��<70�<�d�<:��<T��<`��<Z��<�d�<
0�<���<���<�t�<�<�<h�<���<���<���<���<~��<`   `   ��<���<���<�<��<70�<_H�<�\�<k�<�n�<�j�<�\�<�H�<70�<��<�<���<���<��<d��<���<p��<���<d��<`   `   ���<��<���<���<�r�<�d�<�\�<�Y�<_W�<�W�<�Y�<�\�<�d�<s�<���<x��<��<���<|��<I�<��<��<G�<���<`   `   d��<<��<�9�<F��<߸�<:��<k�<_W�<wP�<_W�<$k�<:��<���<F��<�9�<<��<*��<:�<9W�<~�<P��<~�<W�<:�<`   `   ���<�.�<���<C�<���<T��<�n�<�W�<_W�<vn�<`��<���< C�<{��<�.�<ή�<N)�<��<��<��<��<4��<��<))�<`   `   �Y�<���<, �<2m�<���<`��<�j�<�Y�<$k�<`��<I��<2m�<I �<���<�Y�<
�<���<�!�<�s�<��<�s�<�!�<���<
�<`   `   :��<��<��<&m�<���<Z��<�\�<�\�<:��<���<2m�<|�<!��<O��<­�<��<�6�<Q��<-�<P�<f��<�6�<��<ޭ�<`   `   ���<!��</ �< C�<���<�d�<�H�<�d�<���< C�<I �<!��<���<���<��<���<��<j<�<g�<j<�<��<���<j�<���<`   `   :��<��<���<g��<�r�<
0�<70�<s�<F��<{��<���<O��<���<1=�<=i�<�f�<��<W��<4��<��<g�<Yi�<0=�<���<`   `   Z�<�.�<�9�<���<�<���<��<���<�9�<�.�<�Y�<­�<��<=i�<A��<��<h5�<�k�<�5�<��<��<=i�<��<­�<`   `   ���<\��<���<��<e��<���<�<x��<<��<ή�<
�<��<���<�f�<��<�t�<���<���<ot�<:��<g�<���<��<
�<`   `   ��<��<���<�t�<�J�<�t�<���<��<+��<N)�<���<�6�<��<��<h5�<���<�%�<���<n5�<��<��<�6�<���<N)�<`   `   ���<i��<�<�<���<���<�<�<���<���<:�<��<�!�<Q��<j<�<W��<�k�<���<���<l�<4��<`<�<f��<�!�<��<[�<`   `   S��<h�<���<�b�<��<h�<��<|��<9W�<��<�s�<-�<g�<4��<�5�<ot�<n5�<4��<4g�<-�<�s�<��<W�<|��<`   `   ���<�D�<��<���<�D�<���<d��<I�<~�<��<��<P�<j<�<��<��<:��<��<`<�<-�<��<��<;~�<G�<7��<`   `   K�<#��<�l�<#��<f�<���<���<��<P��<��<�s�<f��<��<g�<��<g�<��<f��<�s�<��<��<��<���<���<`   `   �V�<1
�<W
�<�V�<Z��<���<p��<��<~�<4��<�!�<�6�<���<Yi�<=i�<���<�6�<�!�<��<;~�<��<C��<���<���<`   `   ��<$��<���<�6�<���<���<���<G�<W�<��<���<��<j�<0=�<��<��<���<��<W�<G�<���<���<���<�6�<`   `   Ly�<ay�<]��<�6�<Z��<~��<d��<���<:�<))�<
�<ޭ�<���<���<­�<
�<N)�<[�<|��<7��<���<���<�6�<7��<`   `   ���<���<��<K��<I�<\��<�t�<�4�<��<S��<r�<a]�<y�<a]�<��<S��<���<�4�<�t�<\��<�<K��<��<���<`   `   ���<���<bJ�<��<!;�<z��<,x�<�<O��<b-�<k��<���<���<]��<J-�<p��<;�<�w�<\��<P;�<&��<<J�<���<���<`   `   ��<bJ�<_��<���<\q�<��<;�<� �<�s�<U��<�<��<�<U��<�s�<� �<G�<��<Kq�<���<t��<bJ�<{�<��<`   `   K��<��<���<�P�<��<��<���<��<&<�<�v�<t��<f��<�v�<G<�<��<���<��<��<�P�<���<&��<a��<�l�<�l�<`   `   I�<!;�<\q�<��<���<4K�<3��<Y��<��<�-�<G8�<�-�<f�<Y��<x��<4K�<r��<��<�q�<!;�<"�<+��<���<+��<`   `   \��<z��<��<��<4K�<�y�<���<#��<!��<#��<1��<A��<*��<m��<�y�<dK�<��<���<\��<q��<*��<&��<'��<��<`   `   �t�<,x�<;�<���<3��<���<��<Z��<���<���<���<Z��<��<���<��<���<A�<,x�<�t�<�r�<Ds�<�r�<Us�<�r�<`   `   �4�<�<� �<��<Y��<#��<Z��<W��<���<���<d��<-��<*��<���<��<� �<;�<�4�<�K�<�\�<Af�</f�<�\�<�K�<`   `   ��<O��<�s�<&<�<��<!��<���<���<Ĵ�<���<��<!��<X�<&<�<5t�<O��<���<�"�<�N�<3k�<�t�<3k�<�N�<�"�<`   `   R��<b-�<U��<�v�<�-�<#��<���<���<���<���<1��<�-�<�v�<.��<J-�<h��<���<�6�<�o�<���<ӌ�<�o�<�6�<���<`   `   r�<k��<�<t��<G8�<1��<���<d��<��<1��<
8�<t��<%�<k��<t�<=��<�<`�<���<���<O��<`�<#�<=��<`   `   a]�<���<��<f��<�-�<A��<Z��<-��<!��<�-�<t��<\�<���<w]�<��<ˤ�<�)�<i��<���<Ľ�<{��<�)�<ˤ�<��<`   `   y�<���<�<�v�<f�<*��<��<*��<X�<�v�<%�<���<�x�<:E�<N�<���<�F�<���<B��<���<�F�<���<5�<:E�<`   `   a]�<]��<U��<G<�<Y��<m��<���<���<&<�<.��<k��<w]�<:E�<�.�<��<���<�B�<���<���<�B�<���<��<�.�<3E�<`   `   ��<J-�<�s�<��<x��<�y�<��<��<5t�<J-�<t�<��<N�<��<���<̘�<�	�<�0�<�	�<̘�<���<��<T�<��<`   `   S��<p��<� �<���<4K�<dK�<���<� �<O��<h��<=��<ˤ�<���<���<̘�<�6�<��<���<�6�<��<���<y��<ˤ�</��<`   `   ���<;�<G�<��<r��<��<A�<;�<���<���<�<�)�<�F�<�B�<�	�<��<2��<��<�	�<�B�<�F�<�)�<�<���<`   `   �4�<�w�<��<��<��<���<,x�<�4�<�"�<�6�<`�<i��<���<���<�0�<���<��<�0�<���<���<{��<`�<�6�<#�<`   `   �t�<\��<Kq�<�P�<�q�<\��<�t�<�K�<�N�<�o�<���<���<B��<���<�	�<�6�<�	�<���<g��<���<{��<�o�<�N�<�K�<`   `   \��<P;�<���<���<!;�<q��<�r�<�\�<3k�<���<���<Ľ�<���<�B�<̘�<��<�B�<���<���<���<ӌ�<Tk�<�\�<�r�<`   `   �<&��<t��<&��<"�<*��<Ds�<Af�<�t�<ӌ�<O��<{��<�F�<���<���<���<�F�<{��<{��<ӌ�<rt�<Af�<ps�<*��<`   `   K��<<J�<bJ�<a��<+��<&��<�r�</f�<3k�<�o�<`�<�)�<���<��<��<y��<�)�<`�<�o�<Tk�<Af�<�r�<'��<Z��<`   `   ��<���<{�<�l�<���<'��<Us�<�\�<�N�<�6�<#�<̤�<5�<�.�<T�<̤�<�<�6�<�N�<�\�<ps�<'��<���<�l�<`   `   ���<���<��<�l�<+��<��<�r�<�K�<�"�<���<=��<��<:E�<3E�<��</��<���<#�<�K�<�r�<*��<Z��<�l�<��<`   `   ���<���<7�<�g�<���<�R�<���<�n�<���<(p�<-��<	�<�<	�<N��<(p�<|��<�n�<.��<�R�<~��<�g�<X�<���<`   `   ���<E�<�:�<���<W��<�f�<���<AZ�</��<�&�<i�<���<���<i�<�&�<M��<\Z�<���<xf�<���<���<y:�<G�<���<`   `   7�<�:�<gt�<p��<U�<�~�<e��<�F�<���<x��<@	�<��<I	�<x��<���<�F�<s��<�~�<D�<p��<|t�<�:�< �<�
�<`   `   �g�<���<p��<D�<�L�<���<~��<4�<jp�<]��<���<t��<b��<�p�<�3�<U��<��<
M�<+�<M��<���<�g�<�U�<�U�<`   `   ���<W��<U�<�L�<_��<=��<��<�#�<4J�<�b�<�j�<�b�<J�<�#�<���<=��<��<�L�<��<W��<���<y��<��<y��<`   `   �R�<�f�<�~�<���<=��<���<���<"�<�+�<X5�<e5�<�+�<&�<���<���<h��<��<�~�<xf�<�R�<�E�<'?�<)?�<�E�<`   `   ���<���<e��<~��<��<���<�<c�<��<�<��<c�<+�<���<g��<~��<m��<���<���<@��<���<5��<���<@��<`   `   �n�<AZ�<�F�<4�<�#�<"�<c�<��<!�<@�<��<:�<&�<�#�<�3�<aF�<\Z�<�n�<���<܍�<��<Ք�<ލ�<ր�<`   `   ���</��<���<jp�<4J�<�+�<��<!�<��<!�<��<�+�<J�<jp�<��</��<���< !�<QA�<�V�<�^�<�V�<5A�< !�<`   `   (p�<�&�<x��<]��<�b�<X5�<�<@�<!�<��<e5�<+c�<b��<U��<�&�<=p�<���<���<F�<�-�<�-�<_�<���<ٳ�<`   `   -��<i�<@	�<���<�j�<e5�<��<��<��<e5�<�j�<���<_	�<i�<,��<�.�<ۄ�<`��<���<d�<s��<`��<��<�.�<`   `   	�<���<��<t��<�b�<�+�<c�<:�<�+�<*c�<���<��<���<.	�<��<@��<p[�<���<|��<���<���<U[�<B��<&��<`   `   �<���<I	�<b��<J�<&�<+�<&�<J�<b��<_	�<���<��<j��<E�<-��<�)�<�i�<��<�i�<�)�<-��<E�<j��<`   `   	�<i�<x��<�p�<�#�<���<���<�#�<jp�<U��<i�<.	�<j��<�^�<���<p��<S��<\�<C�<8��<~��<���<�^�<f��<`   `   N��<�&�<���<�3�<���<���<g��<�3�<��<�&�<,��<��<E�<���<��<�<�m�<)��<�m�<�<]��<���<E�<��<`   `   (p�<M��<�F�<U��<=��<h��<~��<aF�</��<=p�<�.�<@��<-��<p��<�<Q��<���<w��<8��<%�<~��<(��<B��<�.�<`   `   |��<\Z�<s��<��<��<��<m��<\Z�<���<���<ۄ�<p[�<�)�<S��<�m�<���<L��<���<�m�<S��<�)�<p[�<��<���<`   `   �n�<���<�~�<
M�<�L�<�~�<���<�n�< !�<���<`��<���<�i�<\�<)��<w��<���<<��<C�<�i�<���<R��<���<!�<`   `   .��<xf�<D�<+�<��<xf�<���<���<QA�<F�<���<|��<��<C�<�m�<8��<�m�<C�<��<|��<���<F�<0A�<���<`   `   �R�<���<p��<M��<W��<�R�<@��<܍�<�V�<�-�<d�<���<�i�<8��<�<%�<S��<�i�<|��<V�<�-�<�V�<ލ�<��<`   `   ~��<���<|t�<���<���<�E�<���<��<�^�<�-�<s��<���<�)�<~��<]��<~��<�)�<���<���<�-�<o^�<��<���<�E�<`   `   �g�<y:�<�:�<�g�<y��<'?�<5��<Ք�<�V�<_�<`��<U[�<-��<���<���<(��<p[�<R��<F�<�V�<��<��<)?�<���<`   `   X�<G�< �<�U�<��<)?�<���<ލ�<5A�<���<��<B��<E�<�^�<E�<B��<��<���<0A�<ލ�<���<)?�<ӹ�<�U�<`   `   ���<���<�
�<�U�<y��<�E�<@��<ր�< !�<ٳ�<�.�<&��<j��<f��<��<�.�<���<!�<���<��<�E�<���<�U�<�
�<`   `   1��<D��<B��<��<�a�<���<s+�<0��<y��<EV�<���<���<��<���<ӛ�<EV�<J��<0��<�+�<���<�a�<��<^��<D��<`   `   D��<��<��<H,�<5y�<���<�,�< ��<���<c�<�P�<j�<	j�<�P�<T�<��<5��<�,�<���<Yy�<S,�<���<��<U��<`   `   B��<��<S�<dS�<]��<���<�/�<�w�<��<x��<1�<��<:�<x��<��<�w�<�/�<���<M��<dS�<e�<��<.��<���<`   `   ��<H,�<dS�<r��<��<W��<�2�<�h�<��<��<F��<:��<��<��<�h�<~2�<l��<0��<^��<FS�<S,�<�<@�<>�<`   `   �a�<5y�<]��<��<���<�<	8�<�\�<�w�<��<P��<��<w�<�\�<;8�<�<u��<��<���<5y�<�a�<�S�<�N�<�S�<`   `   ���<���<���<W��<�<2(�<�=�<�Q�<_�<�f�<�f�<_�<�Q�<�=�<#(�<:�<l��<���<���<���<���<���<���<���<`   `   s+�<�,�<�/�<�2�<	8�<�=�<D�<}I�<{M�<�N�<UM�<}I�<6D�<�=�<�7�<�2�<�/�<�,�<u+�<v+�<�+�<f+�<�+�<v+�<`   `   0��< ��<�w�<�h�<�\�<�Q�<}I�<jE�<�B�<�B�<vE�<ZI�<�Q�<�\�<�h�<�w�<5��<A��<l��<���<���<���<���<���<`   `   y��<���<��<��<�w�<_�<{M�<�B�<�=�<�B�<�M�<_�<uw�<��<D��<���<R��<)�<;4�<�C�<cI�<�C�<%4�<)�<`   `   EV�<c�<x��<��<��<�f�<�N�<�B�<�B�<fN�<�f�<;��<��<Z��<T�<WV�<ӈ�<޳�<P��<X��<b��<d��<��<���<`   `   ���<�P�<1�<F��<P��<�f�<UM�<vE�<�M�<�f�< ��<F��<L�<�P�<���<Y��<�"�<+T�<�s�<�~�<�s�<+T�<�"�<Y��<`   `   ���<j�<��<:��<��<_�<}I�<ZI�<_�<;��<F��<q�<	j�<���<O$�<Jy�<��<2��<�<�<=��<Կ�<My�<^$�<`   `   ��<	j�<:�<��<w�<�Q�<6D�<�Q�<uw�<��<L�<	j�<���<�E�<l��<��<�V�<K��<֔�<K��<�V�<��<Z��<�E�<`   `   ���<�P�<x��<��<�\�<�=�<�=�<�\�<��<Z��<�P�<���<�E�<���<�5�<m��<e��<g��<S��<O��<x��<�5�<���<�E�<`   `   ӛ�<T�<��<�h�<;8�<#(�<�7�<�h�<D��<T�<���<O$�<l��<�5�<��<'�<.A�</U�<WA�<'�<ת�<�5�<l��<O$�<`   `   EV�<��<�w�<~2�<�<:�<�2�<�w�<���<WV�<Y��<Jy�<��<m��<'�<rX�<���<l��<_X�<6�<x��<��<My�<M��<`   `   J��<5��<�/�<l��<u��<l��<�/�<5��<R��<ӈ�<�"�<��<�V�<e��<.A�<���<���<���<2A�<e��<�V�<��<�"�<ӈ�<`   `   0��<�,�<���<0��<��<���<�,�<A��<)�<޳�<+T�<2��<K��<g��</U�<l��<���<>U�<S��<H��<=��<T�<��<C�<`   `   �+�<���<M��<^��<���<���<u+�<l��<;4�<P��<�s�<�<֔�<S��<WA�<_X�<2A�<S��<��<�<�s�<P��<4�<l��<`   `   ���<Yy�<dS�<FS�<5y�<���<v+�<���<�C�<X��<�~�<�<K��<O��<'�<6�<e��<H��<�<�~�<b��<�C�<���<T+�<`   `   �a�<S,�<e�<S,�<�a�<���<�+�<���<cI�<b��<�s�<=��<�V�<x��<ت�<x��<�V�<=��<�s�<b��<>I�<���<,�<���<`   `   ��<���<��<�<�S�<���<f+�<���<�C�<d��<+T�<Կ�<��<�5�<�5�<��<��<T�<P��<�C�<���<D+�<���<�S�<`   `   ^��<��<.��<@�<�N�<���<�+�<���<%4�<��<�"�<My�<Z��<���<l��<My�<�"�<��<4�<���<,�<���<[N�<@�<`   `   D��<U��<���<>�<�S�<���<v+�<���<)�<���<Y��<^$�<�E�<�E�<O$�<M��<ӈ�<C�<l��<T+�<���<�S�<@�<p��<`   `   �7�<>B�<~_�<��<���<��<�b�<Բ�<d��<�@�<�s�<7��<���<7��<�s�<�@�<B��<Բ�<�b�<��<���<��<�_�<>B�<`   `   >B�<�R�<�s�<���<a��<?�<�b�<���<���<��<�;�<�N�<�N�<�;�<��<���<���<�b�<1�<|��<���<rs�<�R�<KB�<`   `   }_�<�s�<��<`��<{��<�+�<�d�<���<���<r��<��<��<��<r��<���<���<�d�<�+�<n��<`��< ��<�s�<n_�<{X�<`   `   ��<���<`��<���<��<�;�<&g�<*��<1��<���<��<���<���<E��<��<g�<�;�<��<���<J��<���<!��<3��<1��<`   `   ���<a��<{��<��<N-�<�L�<sj�<ф�<��<6��<���<6��<ܘ�<ф�<�j�<�L�<$-�<��<���<a��<���<���<��<���<`   `   ��<?�<�+�<�;�<�L�<a^�<�n�<0|�<?��<I��<R��<R��<2|�<�n�<W^�<�L�<�;�<�+�<1�<��<��<��<��<��<`   `   �b�<�b�<�d�<&g�<sj�<�n�<Lr�<>u�<�w�<�w�<�w�<>u�<dr�<�n�<cj�<&g�<�d�<�b�<�b�<b�<>b�<Ob�<Cb�<b�<`   `   Բ�<���<���<*��<ф�<0|�<>u�<|q�<o�<o�<�q�<%u�<2|�<��<��<z��<���<��<Լ�<L��<1��<)��<N��<��<`   `   d��<���<���<1��<��<?��<�w�<o�<�k�<o�<�w�<?��<՘�<1��<��<���<H��<��<�'�<�3�<K7�<�3�<�'�<��<`   `   �@�<��<r��<���<6��<I��<�w�<o�<o�<�w�<R��<Q��<���<\��<��<�@�<!f�<���<���<;��<C��<���<���<f�<`   `   �s�<�;�<��<��<���<R��<�w�<�q�<�w�<R��<���<��<��<�;�<�s�<#��<���<^��<��<��<��<^��<��<#��<`   `   7��<�N�<��<���<6��<R��<>u�<%u�<?��<Q��<��<��<�N�<D��<���<P�<�K�<�p�<���<���<q�<zK�<R�<���<`   `   ���<�N�<��<���<ܘ�<2|�<dr�<2|�<՘�<���<��<�N�<���<���<�?�<4��<s��<!��<p��<!��<{��<4��<x?�<���<`   `   7��<�;�<r��<E��<ф�<�n�<�n�<��<1��<\��<�;�<D��<���<xM�<á�<��<��<<3�<.3�<��<$��<͡�<{M�<���<`   `   �s�<��<���<��<�j�<W^�<cj�<��<��<��<�s�<���<�?�<á�<���<|9�<c�<�q�<�c�<|9�<���<á�<�?�<���<`   `   �@�<���<���<g�<�L�<�L�<&g�<z��<���<�@�<#��<P�<4��<��<|9�<ht�<���<���<Zt�<�9�<$��<2��<R�<��<`   `   B��<���<�d�<�;�<$-�<�;�<�d�<���<H��<!f�<���<�K�<s��<��<c�<���<c��<���<�c�<��<m��<�K�<��<!f�<`   `   Բ�<�b�<�+�<��<��<�+�<�b�<��<��<���<^��<�p�<!��<<3�<�q�<���<���< r�<.3�<��<q�<T��<���<��<`   `   �b�<1�<n��<���<���<1�<�b�<Լ�<�'�<���<��<���<p��<.3�<�c�<Zt�<�c�<.3�<���<���<��<���<�'�<Լ�<`   `   ��<|��<`��<J��<a��<��<b�<L��<�3�<;��<��<���<!��<��<|9�<�9�<��<��<���<��<C��<�3�<N��<�a�<`   `   ���<���< ��<���<���<��<>b�<1��<K7�<C��<��<q�<{��<$��<���<$��<m��<q�<��<C��<07�<1��<Ub�<��<`   `   ��<rs�<�s�<!��<���<��<Ob�<)��<�3�<���<^��<zK�<4��<͡�<á�<2��<�K�<T��<���<�3�<1��<5b�<��<���<`   `   �_�<�R�<n_�<3��<��<��<Cb�<N��<�'�<���<��<R�<x?�<{M�<�?�<R�<��<���<�'�<N��<Ub�<��<Ѽ�<3��<`   `   >B�<KB�<{X�<1��<���<��<b�<��<��<f�<#��<���<���<���<���<��<!f�<��<Լ�<�a�<��<���<3��<eX�<`   `   ���<a��<G��<��<\�<�N�<���<���<���<�.�<�T�<�l�<�t�<�l�<�T�<�.�<���<���<���<�N�<H�<��<S��<a��<`   `   a��<V��<���<���<�%�<�V�<"��<���<���<H�<�*�<�8�<�8�<�*�<B�<���<���<��<�V�<�%�<���<���<X��<i��<`   `   G��<���<���<��<�6�<z`�<9��<H��<��<	��<V�<��<Z�<	��<��<H��<?��<z`�<�6�<��<���<���<>��<���<`   `   ��<���<��<�+�<�J�<(l�<��<2��<@��<���<���<���<���<K��<,��<��<1l�<�J�<�+�<��<���<��<��<��<`   `   \�<�%�<�6�<�J�<Sa�<y�<���<&��<���<���<���<���<���<&��<���<y�<:a�<�J�<�6�<�%�<P�<F�<j�<F�<`   `   �N�<�V�<z`�<(l�<y�<(��<��<���<f��<ͥ�<ҥ�<q��<���<Ӑ�<"��<y�<1l�<m`�<�V�<�N�<pI�<sF�<uF�<lI�<`   `   ���<"��<9��<��<���<��<:��<���<0��<З�<��<���<H��<��<���<��<=��<"��<���<k��<���<j��<���<k��<`   `   ���<���<H��<2��<&��<���<���<���<s��<~��<���<���<���<5��<,��<;��<���<���<���<~��<p��<l��<��<���<`   `   ���<���<��<@��<���<f��<0��<s��<`��<s��<9��<f��<���<@��</��<���<���<��< �<�$�<�'�<�$�<��<��<`   `   �.�<H�<	��<���<���<ͥ�<З�<~��<s��<���<ҥ�<���<���<���<B�</�<�J�<�a�<�r�<k{�<p{�<�r�<�a�<�J�<`   `   �T�<�*�<V�<���<���<ҥ�<��<���<9��<ҥ�<���<���<a�<�*�<�T�<\|�<ڞ�<L��<|��<j��<o��<L��<��<\|�<`   `   �l�<�8�<��<���<���<q��<���<���<f��<���<���<��<�8�<�l�<B��<���<���<��<1�<9�<��<���<���<I��<`   `   �t�<�8�<Z�<���<���<���<H��<���<���<���<a�<�8�<�t�<���<���<@�<LD�<�\�<)e�<�\�<PD�<@�<���<���<`   `   �l�<�*�<	��<K��<&��<Ӑ�<��<5��<@��<���<�*�<�l�<���<F��<3�<�e�<S��<���<���<J��<�e�<3�<G��<���<`   `   �T�<B�<��<,��<���<"��<���<,��</��<B�<�T�<B��<���<3�<�q�<��<���<h��<���<��<�q�<3�<���<B��<`   `   �.�<���<H��<��<y�<y�<��<;��<���</�<\|�<���<@�<�e�<��<���<��<��<���<��<�e�<?�<���<V|�<`   `   ���<���<?��<1l�<:a�<1l�<=��<���<���<�J�<ڞ�<���<LD�<S��<���<��<0��<��<���<S��<HD�<���<ޞ�<�J�<`   `   ���<��<z`�<�J�<�J�<m`�<"��<���<��<�a�<L��<��<�\�<���<h��<��<��<n��<���<�\�<��<G��<�a�<��<`   `   ���<�V�<�6�<�+�<�6�<�V�<���<���< �<�r�<|��<1�<)e�<���<���<���<���<���<2e�<1�<}��<�r�<��<���<`   `   �N�<�%�<��<��<�%�<�N�<k��<~��<�$�<k{�<j��<9�<�\�<J��<��<��<S��<�\�<1�<e��<p{�<�$�<��<\��<`   `   H�<���<���<���<P�<pI�<���<p��<�'�<p{�<o��<��<PD�<�e�<�q�<�e�<HD�<��<}��<p{�<�'�<p��<É�<pI�<`   `   ��<���<���<��<F�<sF�<j��<l��<�$�<�r�<L��<���<@�<3�<3�<?�<���<G��<�r�<�$�<p��<[��<uF�<U�<`   `   S��<X��<>��<��<j�<uF�<���<��<��<�a�<��<���<���<G��<���<���<ޞ�<�a�<��<��<É�<uF�<Y�<��<`   `   a��<i��<���<��<F�<lI�<k��<���<��<�J�<\|�<I��<���<���<B��<V|�<�J�<��<���<\��<pI�<U�<��<���<`   `   F��<Y�<y�<.�<�P�<�x�<ڤ�<���<q��<~�<�;�<�M�<)S�<�M�<�;�<~�<k��<���<��<�x�<�P�<.�<|�<Y�<`   `   Y�<��<j�<�9�<�Z�<�~�<���<8��<���<,	�<g�<�'�<�'�<f�<*	�< ��<;��<���<�~�<�Z�<:�<g�<��<[�<`   `   y�<j�<(2�<{J�<vg�<���<=��<���<���<���<n��<�<n��<���<���<���<>��<���<ug�<{J�<)2�<j�<x�<��<`   `   .�<�9�<{J�<F_�<�v�<��<���<a��<c��<���<���<���<���<e��<_��<���<��<�v�<D_�<xJ�<:�<.�<X(�<X(�<`   `   �P�<�Z�<vg�<�v�<��<`��<ƨ�<���<���<���<@��<���<���<���<̨�<`��<���<�v�<|g�<�Z�<�P�<�J�<H�<�J�<`   `   �x�<�~�<���<��<`��<j��<P��<2��<��<��<��<��<3��<M��<g��<d��<��<���<�~�<�x�<Fu�<�r�<�r�<Du�<`   `   ڤ�<���<=��<���<ƨ�<P��<���<��<��<���<��<��<���<P��<Ĩ�<���<=��<���<ۤ�<A��<W��<+��<Y��<A��<`   `   ���<8��<���<a��<���<2��<��<��<���<���<��<��<3��<���<_��<���<;��<���<���<~��<x��<v��<~��<���<`   `   q��<���<���<c��<���<��<��<���<���<���<��<��<���<c��<���<���<l��<��<��<��<��<��<��<��<`   `   ~�<,	�<���<���<���<��<���<���<���<���<��<���<���<���<*	�<��<�4�<6F�<�R�<�X�<�X�<�R�<6F�<�4�<`   `   �;�<g�<n��<���<@��<��<��<��<��<��<;��<���<p��<g�<�;�<�X�<�r�<u��<���<���<���<u��<�r�<�X�<`   `   �M�<�'�<�<���<���<��<��<��<��<���<���<�<�'�<�M�<>s�<9��<9��<l��<���<���<m��<6��<9��<@s�<`   `   )S�<�'�<n��<���<���<3��<���<3��<���<���<p��<�'�<'S�<T��<Z��<���<���<���<��<���<���<���<X��<T��<`   `   �M�<f�<���<e��<���<M��<P��<���<c��<���<g�<�M�<T��<���<���<�<��<H-�<E-�<��<�<���<���<S��<`   `   �;�<*	�<���<_��<̨�<g��<Ĩ�<_��<���<*	�<�;�<>s�<Z��<���<G�<�0�<2G�<�N�<8G�<�0�<C�<���<[��<>s�<`   `   ~�< ��<���<���<`��<d��<���<���<���<��<�X�<9��<���<�<�0�<\P�<Y`�<V`�<ZP�<�0�<�<���<9��<�X�<`   `   k��<;��<>��<��<���<��<=��<;��<l��<�4�<�r�<9��<���<��<2G�<Y`�<�h�<Y`�<3G�<��<���<9��<�r�<�4�<`   `   ���<���<���<�v�<�v�<���<���<���<��<6F�<u��<l��<���<H-�<�N�<V`�<Y`�<�N�<E-�<���<m��<t��<6F�<��<`   `   ��<�~�<ug�<D_�<|g�<�~�<ۤ�<���<��<�R�<���<���<��<E-�<8G�<ZP�<3G�<E-�<��<���<���<�R�<��<���<`   `   �x�<�Z�<{J�<xJ�<�Z�<�x�<A��<~��<��<�X�<���<���<���<��<�0�<�0�<��<���<���<���<�X�<��<~��<=��<`   `   �P�<:�<)2�<:�<�P�<Fu�<W��<x��<��<�X�<���<m��<���<�<C�<�<���<m��<���<�X�<��<x��<[��<Fu�<`   `   .�<g�<j�<.�<�J�<�r�<+��<v��<��<�R�<u��<6��<���<���<���<���<9��<t��<�R�<��<x��<'��<�r�<�J�<`   `   |�<��<x�<X(�<H�<�r�<Y��<~��<��<6F�<�r�<9��<X��<���<[��<9��<�r�<6F�<��<~��<[��<�r�<{H�<X(�<`   `   Y�<[�<��<X(�<�J�<Du�<A��<���<��<�4�<�X�<@s�<T��<S��<>s�<�X�<�4�<��<���<=��<Fu�<�J�<X(�<��<`   `   ;�<�?�<L�<�_�<`y�<��<!��<N��<���<��<(�<Z5�<�9�<Z5�<(�<��<���<N��<��<��<iy�<�_�<L�<�?�<`   `   �?�<G�<�T�<jh�<ɀ�<V��<��<���<��<��<V�<��<��<Y�<��<��<���<���<Y��<���<ih�<�T�<G�<�?�<`   `   L�<�T�<pb�<�t�<\��<���<���<���<���<���<b��<���<^��<���<���<���<���<���<`��<�t�<kb�<�T�<L�<	I�<`   `   �_�<jh�<�t�<G��<���<��<߹�<���<=��<���<���<���<���<8��<���<��<��<���<J��<�t�<ih�<�_�<4[�<6[�<`   `   `y�<ɀ�<\��<���<<��<׮�<���<���<)��<S��<c��<S��</��<���<���<׮�<G��<���<R��<ɀ�<ey�<�t�<bs�<�t�<`   `   ��<V��<���<��<׮�<���<���<���<���<��<|��<���<���<���<���<Ю�<��<���<Y��<��<���<S��<Q��<���<`   `   !��<��<���<߹�<���<���<C��<ؽ�<0��<���<8��<ؽ�<<��<���<���<߹�<���<��<"��<���<M��<���<N��<���<`   `   N��<���<���<���<���<���<ؽ�<}��<��<��<z��<߽�<���<���<���<���<���<J��<��<���<���<���<���<��<`   `   ���<��<���<=��<)��<���</��<��<9��<��<+��<���<1��<=��<���<��<���<�<@	�<,�<�<,�<D	�<�<`   `   ��<��<���<���<S��<��<���<��<��<��<|��<K��<���<���<��<��<�#�<{/�<�8�<�=�<�=�<�8�<z/�<�#�<`   `   (�<V�<b��<���<c��<|��<8��<z��<+��<|��<n��<���<[��<V�<(�<4>�<�P�<Z_�<�h�<�k�<�h�<Z_�<�P�<4>�<`   `   Z5�<��<���<���<S��<���<ؽ�<߽�<���<K��<���<���<��<U5�<CQ�<oj�<D�<���<���<���<��<G�<nj�<AQ�<`   `   �9�<��<^��<���</��<���<<��<���<1��<���<[��<��<�9�<N[�<�z�<���<���<·�<���<·�<���<���<�z�<N[�<`   `   Z5�<Y�<���<8��<���<���<���<���<=��<���<V�<U5�<N[�<��<\��<���<O��<���<���<R��<���<Z��<��<M[�<`   `   (�<��<���<���<���<���<���<���<���<��<(�<CQ�<�z�<\��<D��<���<���<g��<���<���<G��<\��<�z�<CQ�<`   `   ��<��<���<��<׮�<Ю�<߹�<���<��<��<4>�<oj�<���<���<���<���<���<���<���<���<���<���<nj�<7>�<`   `   ���<���<���<��<G��<��<���<���<���<�#�<�P�<D�<���<O��<���<���<��<���<���<O��<���<D�<�P�<�#�<`   `   N��<���<���<���<���<���<��<J��<�<{/�<Z_�<���<·�<���<g��<���<���<e��<���<·�<��<]_�<z/�<��<`   `   ��<Y��<`��<J��<R��<Y��<"��<��<@	�<�8�<�h�<���<���<���<���<���<���<���<���<���<�h�<�8�<G	�<��<`   `   ��<���<�t�<�t�<ɀ�<��<���<���<,�<�=�<�k�<���<·�<R��<���<���<O��<·�<���<�k�<�=�<'�<���<Ǹ�<`   `   iy�<ih�<kb�<ih�<ey�<���<M��<���<�<�=�<�h�<��<���<���<G��<���<���<��<�h�<�=�<$�<���<G��<���<`   `   �_�<�T�<�T�<�_�<�t�<S��<���<���<,�<�8�<Z_�<G�<���<Z��<\��<���<D�<]_�<�8�<'�<���< ��<Q��<�t�<`   `   L�<G�<L�<4[�<bs�<Q��<N��<���<D	�<z/�<�P�<nj�<�z�<��<�z�<nj�<�P�<z/�<G	�<���<G��<Q��<ks�<4[�<`   `   �?�<�?�<	I�<6[�<�t�<���<���<��<�<�#�<4>�<AQ�<N[�<M[�<CQ�<7>�<�#�<��<��<Ǹ�<���<�t�<4[�<I�<`   `   bh�<�k�<�t�<~��<��<2��<���<M��<���<J	�<��<]"�<�%�<]"�<��<J	�<���<M��<���<2��<��<~��<�t�<�k�<`   `   �k�<q�<A{�<��<��<���<���<d��<���<j��<a�<R�<R�<h�<p��<���<\��<���<���<��<��<P{�<q�<�k�<`   `   �t�<A{�<���<y��<���<���<���<���<���<7��<���<P��<���<7��<���<���<���<���<���<y��<���<A{�<�t�<zr�<`   `   ~��<��<y��<
��<��<��<J��<���<x��<���<��<��<���<k��<���<[��<v��<���<��<���<��<u��<��<��<`   `   ��<��<���<��<���<\��<m��<���<��<\��<n��<\��<��<���<V��<\��<��<��<���<��< ��<��<��<��<`   `   2��<���<���<��<\��<y��<<��<���<���<���<���<|��<���<M��<��<J��<v��<���<���<)��<D��< ��<���<H��<`   `   ���<���<���<J��<m��<<��<���<���<`��<���<t��<���<���<<��<y��<J��<���<���<���<���<v��<���<u��<���<`   `   M��<d��<���<���<���<���<���<���<p��<c��<���<���<���<{��<���<���<\��<D��<���<���<���<���<���<~��<`   `   ���<���<���<x��<��<���<`��<p��<���<p��<V��<���<��<x��<���<���<���<���<M�<��<V�<��<W�<���<`   `   J	�<j��<7��<���<\��<���<���<c��<p��<���<���<J��<���<F��<p��<@	�<��<�<%�<L(�<H(�<%�<�<��<`   `   ��<a�<���<��<n��<���<t��<���<V��<���<���<��<���<a�<��<�(�<g6�<�A�<LH�<�J�<XH�<�A�<`6�<�(�<`   `   ]"�<R�<P��<��<\��<|��<���<���<���<J��<��<_��<R�<T"�<7�<eI�<Y�<�c�<<i�<4i�<�c�<Y�<cI�<�6�<`   `   �%�<R�<���<���<��<���<���<���<��<���<���<R�<�%�<K>�<U�<9i�<�x�<V��<��<V��<�x�<9i�<U�<K>�<`   `   ]"�<h�<7��<k��<���<M��<<��<{��<x��<F��<a�<T"�<K>�<EY�<�q�<;��<���<���<���<���<7��<�q�<BY�<K>�<`   `   ��<p��<���<���<V��<��<y��<���<���<p��<��<7�<U�<�q�<Ȋ�<���<ȩ�<���<���<���<ъ�<�q�<U�<7�<`   `   J	�<���<���<[��<\��<J��<J��<���<���<@	�<�(�<eI�<9i�<;��<���<V��<8��<@��<^��<���<7��<9i�<cI�<�(�<`   `   ���<\��<���<v��<��<v��<���<\��<���<��<g6�<Y�<�x�<���<ȩ�<8��<˻�<8��<Ʃ�<���<�x�<Y�<b6�<��<`   `   M��<���<���<���<��<���<���<D��<���<�<�A�<�c�<V��<���<���<@��<8��<���<���<V��<�c�<�A�<�<u��<`   `   ���<���<���<��<���<���<���<���<M�<%�<LH�<<i�<��<���<���<^��<Ʃ�<���<��<<i�<IH�<%�<\�<���<`   `   2��<��<y��<���<��<)��<���<���<��<L(�<�J�<4i�<V��<���<���<���<���<V��<<i�<�J�<H(�<��<���<���<`   `   ��<��<���<��< ��<D��<v��<���<V�<H(�<XH�<�c�<�x�<7��<ъ�<7��<�x�<�c�<IH�<H(�<g�<���<h��<D��<`   `   ~��<P{�<A{�<u��<��< ��<���<���<��<%�<�A�<Y�<9i�<�q�<�q�<:i�<Y�<�A�<%�<��<���<���<���<m��<`   `   �t�<q�<�t�<��<��<���<u��<���<W�<�<`6�<cI�<U�<BY�<U�<cI�<b6�<�<\�<���<h��<���<��<��<`   `   �k�<�k�<zr�<��<��<H��<���<~��<���<��<�(�<�6�<K>�<K>�<7�<�(�<��<u��<���<���<D��<m��<��<�r�<`   `   d��<3��<��<��<���<E��<l��<��<��<� �<{�<�<T�<�<h�<� �<,��<��<F��<E��<���<��<��<3��<`   `   3��<���<��<<��<���<��<��<v��<���<b��<S��<f�<e�<\��<l��<���<h��<2��<��<k��<5��</��<���<&��<`   `   ��<��<��<���<��</��<@��<���<���<e��<\��<���<T��<e��<���<���<5��</��<��<���<ܞ�<��<+��<ɐ�<`   `   ��<<��<���<��<V��<_��<��<'��<@��<,��<O��<X��<+��<-��<1��<��<Q��<<��<��<��<5��<��<��<��<`   `   ���<���<��<V��<Z��<���<���<;��<���<��<���<��<���<;��<c��<���<���<V��<��<���<���<��<M��<��<`   `   E��<��</��<_��<���<��<���<���<C��<���<���<0��<���<���<$��<���<Q��<E��<��<8��<��<���<���<��<`   `   l��<��<@��<��<���<���<��<���<���<*��< ��<���<��<���<���<��<8��<��<l��<���<���<Y��<���<���<`   `   ��<v��<���<'��<;��<���<���<���<s��<`��<���<���<���<!��<1��<��<h��<��<���<���<���<���<���<���<`   `   ��<���<���<@��<���<C��<���<s��<V��<s��<���<C��<���<@��<���<���<&��<���<��<u��<l��<u��<&��<���<`   `   � �<b��<e��<,��<��<���<*��<`��<s��<C��<���<��<+��<{��<l��<z �<��<R�<��<��<��<��<O�<��<`   `   {�<S��<\��<O��<���<���< ��<���<���<���<���<O��<G��<S��<�<��<$"�<@*�<�.�<%1�</�<@*�<"�<��<`   `   �<f�<���<X��<��<0��<���<���<C��<��<O��<���<e�<�<m"�<<0�<�;�<YC�<�G�<�G�<RC�<�;�<90�<c"�<`   `   T�<e�<T��<+��<���<���<��<���<���<+��<G��<e�<b�<�'�<*9�<�G�<�R�<wZ�<]�<wZ�<�R�<�G�<69�<�'�<`   `   �<\��<e��<-��<;��<���<���<!��<@��<{��<S��<�<�'�<-<�<+N�<�\�<�g�<�l�<�l�<�g�<�\�<"N�<*<�<�'�<`   `   h�<l��<���<1��<c��<$��<���<1��<���<l��<�<m"�<*9�<+N�<`�<�n�<iw�<�y�<Nw�<�n�<*`�<+N�<+9�<m"�<`   `   � �<���<���<��<���<���<��<��<���<z �<��<<0�<�G�<�\�<�n�<%{�<P��<^��<2{�<n�<�\�<�G�<90�<��<`   `   ,��<h��<5��<Q��<���<Q��<8��<h��<&��<��<$"�<�;�<�R�<�g�<iw�<P��<���<P��<ew�<�g�< S�<�;�<"�<��<`   `   ��<2��</��<<��<V��<E��<��<��<���<R�<@*�<YC�<wZ�<�l�<�y�<^��<P��<�y�<�l�<xZ�<RC�<I*�<O�<���<`   `   F��<��<��<��<��<��<l��<���<��<��<�.�<�G�<]�<�l�<Nw�<2{�<ew�<�l�<�\�<�G�<�.�<��<,��<���<`   `   E��<k��<���<��<���<8��<���<���<u��<��<%1�<�G�<wZ�<�g�<�n�<n�<�g�<xZ�<�G�</1�<��<b��<���<���<`   `   ���<5��<ܞ�<5��<���<��<���<���<l��<��</�<RC�<�R�<�\�<*`�<�\�< S�<RC�<�.�<��<���<���<���<��<`   `   ��</��<��<��<��<���<Y��<���<u��<��<@*�<�;�<�G�<"N�<+N�<�G�<�;�<I*�<��<b��<���<r��<���<˨�<`   `   ��<���<+��<��<M��<���<���<���<&��<O�<"�<90�<69�<*<�<+9�<90�<"�<O�<,��<���<���<���<j��<��<`   `   3��<&��<ɐ�<��<��<��<���<���<���<��<��<c"�<�'�<�'�<m"�<��<��<���<���<���<��<˨�<��<ߐ�<`   `   ���<��<5��<5��<��<���<��<F��<���<��<��<��<	�<��<o�<��<��<F��<���<���<0��<5��<��<��<`   `   ��<P��<���<��<��<���<��<���<���<��<U��<_��<\��<_��<��<���<���<$��<��<��<��<��<M��<ء�<`   `   5��<���<
��<��<#��<���<���<q��<&��<!��<���<��<���<!��</��<q��<���<���<2��<��<���<���<G��<���<`   `   5��<��<��<���<O��<r��<���<���<5��<a��<��<��<^��<��<���<���<_��</��<���<���<��<%��<F��<H��<`   `   ��<��<#��<O��<���<0��<���<���<p��<"��<���<"��<���<���<���<0��<��<O��<���<��< ��<���<���<���<`   `   ���<���<���<r��<0��<���<��<��<\��<"��<��<E��<
��<6��<���<��<_��<���<��<���<��<���<���<!��<`   `   ��<��<���<���<���<��<��<���<Z��<q��<{��<���<���<��<���<���<���<��<��<S��<���<��<���<S��<`   `   F��<���<q��<���<���<��<���<���<���<���<���<���<
��<���<���<���<���<6��<O��<���<��<%��<���<=��<`   `   ���<���<&��<5��<p��<\��<Z��<���<��<���<F��<\��<���<5��<���<���<��<���<#��<���<���<���<7��<���<`   `   ��<��<!��<a��<"��<"��<q��<���<���<���<��<��<^��<;��<��<���<���<��<�<�
�<�
�<��<��<���<`   `   ��<U��<���<��<���<��<{��<���<F��<��<���<��<���<U��<��<�
�<�<��<�<��<��<��<�<�
�<`   `   ��<_��<��<��<"��<E��<���<���<\��<��<��<��<\��<��<��<>�<d$�<�*�<h-�<W-�<�*�<w$�<<�<��<`   `   	�<\��<���<^��<���<
��<���<
��<���<^��<���<\��<%	�<K�<�"�<�-�<�5�<�;�<=�<�;�<�5�<�-�<�"�<K�<`   `   ��<_��<!��<��<���<6��<��<���<5��<;��<U��<��<K�<�$�<!2�<`=�<�D�<�H�<�H�<�D�<V=�<2�<�$�<N�<`   `   o�<��</��<���<���<���<���<���<���<��<��<��<�"�<!2�<�?�<J�<�P�<bS�<}P�<J�<@�<!2�<�"�<��<`   `   ��<���<q��<���<0��<��<���<���<���<���<�
�<>�<�-�<`=�<J�<�R�<�W�<X�<�R�<J�<V=�<�-�<<�<�
�<`   `   ��<���<���<_��<��<_��<���<���<��<���<�<d$�<�5�<�D�<�P�<�W�<�Y�<�W�<�P�<�D�<�5�<d$�<�<���<`   `   F��<$��<���</��<O��<���<��<6��<���<��<��<�*�<�;�<�H�<bS�<X�<�W�<TS�<�H�<�;�<�*�<��<��<���<`   `   ���<��<2��<���<���<��<��<O��<#��<�<�<h-�<=�<�H�<}P�<�R�<�P�<�H�<�<�<h-�<~�<�<<��<O��<`   `   ���<��<��<���<��<���<S��<���<���<�
�<��<W-�<�;�<�D�<J�<J�<�D�<�;�<h-�<��<�
�<���<���<q��<`   `   0��<��<���<��< ��<��<���<��<���<�
�<��<�*�<�5�<V=�<@�<V=�<�5�<�*�<~�<�
�<��<��<���<��<`   `   5��<��<���<%��<���<���<��<%��<���<��<��<w$�<�-�<2�<!2�<�-�<d$�<��<�<���<��</��<���<���<`   `   ��<M��<G��<F��<���<���<���<���<7��<��<�<<�<�"�<�$�<�"�<<�<�<��<<��<���<���<���<շ�<F��<`   `   ��<ء�<���<H��<���<!��<S��<=��<���<���<�
�<��<K�<N�<��<�
�<���<���<O��<q��<��<���<F��<ť�<`   `   ��<α�<µ�<��<8��<��<=��<:��<���<���<���<���<&��<���<���<���<���<:��<��<��<h��<��<���<α�<`   `   α�<��<���<���<���<��<H��<���<2��<$��<���<���<���<���<4��<��<���<i��<1��<���<��<���<��<���<`   `   µ�<���<��<���<0��<t��<��<#��<���<L��<��<���<��<L��<���<#��<���<t��<>��<���<��<���<ӵ�<��<`   `   ��<���<���<r��<���<Y��<p��<3��<��<%��<���<���< ��<���<D��<���<B��<^��<���<���<��<���<`��<a��<`   `   8��<���<0��<���<���<v��<���<t��<��<@��<���<@��<5��<t��<Y��<v��<3��<���<���<���<U��<n��<&��<n��<`   `   ��<��<t��<Y��<v��<���<���<L��<T��</��<%��<;��<G��<��<���<S��<B��<���<1��<��<��<���<���<��<`   `   =��<H��<��<p��<���<���<���<��<��<���<8��<��<���<���<���<p��<���<H��<8��<���<���<Z��<���<���<`   `   :��<���<#��<3��<t��<L��<��<���<���<���<���<2��<G��<Q��<D��<?��<���<)��<���<d��<���<���<c��<���<`   `   ���<2��<���<��<��<T��<��<���<���<���<���<T��<?��<��<���<2��<���<Y��<���<���</��<���<��<Y��<`   `   ���<$��<L��<%��<@��</��<���<���<���<���<%��<��< ��<h��<4��<���<X��<���<���<+��<��<���<���<o��<`   `   ���<���<��<���<���<%��<8��<���<���<%��<���<���<���<���<���<���<��<h	�<O�<��<q�<h	�<��<���<`   `   ���<���<���<���<@��<;��<��<2��<T��<��<���<��<���<���< �<��<��<��<��<l�<��<��<��<�<`   `   &��<���<��< ��<5��<G��<���<G��<?��< ��<���<���<;��<E�<��<��<��<�#�<B%�<�#�<��<��<��<E�<`   `   ���<���<L��<���<t��<��<���<Q��<��<h��<���<���<E�<��<��<i%�<�*�<�-�<�-�<�*�<\%�<��<��<I�<`   `   ���<4��<���<D��<Y��<���<���<D��<���<4��<���< �<��<��<4'�<�.�<�3�<X5�<q3�<�.�<R'�<��<��< �<`   `   ���<��<#��<���<v��<S��<p��<?��<2��<���<���<��<��<i%�<�.�<5�<9�<9�<,5�<�.�<\%�<��<��<���<`   `   ���<���<���<B��<3��<B��<���<���<���<X��<��<��<��<�*�<�3�<9�<v:�<9�<�3�<�*�<��<��<��<X��<`   `   :��<i��<t��<^��<���<���<H��<)��<Y��<���<h	�<��<�#�<�-�<X5�<9�<9�<G5�<�-�<�#�<��<s	�<���<@��<`   `   ��<1��<>��<���<���<1��<8��<���<���<���<O�<��<B%�<�-�<q3�<,5�<�3�<�-�<(%�<��<Q�<���<��<���<`   `   ��<���<���<���<���<��<���<d��<���<+��<��<l�<�#�<�*�<�.�<�.�<�*�<�#�<��<��<��<���<c��<��<`   `   h��<��<��<��<U��<��<���<���</��<��<q�<��<��<\%�<R'�<\%�<��<��<Q�<��<T��<���<t��<��<`   `   ��<���<���<���<n��<���<Z��<���<���<���<h	�<��<��<��<��<��<��<s	�<���<���<���<{��<���<K��<`   `   ���<��<ӵ�<`��<&��<���<���<c��<��<���<��<��<��<��<��<��<��<���<��<c��<t��<���<J��<`��<`   `   α�<���<��<a��<n��<��<���<���<Y��<o��<���<�<E�<I�< �<���<X��<@��<���<��<��<K��<`��<��<`   `   ��<޼�<���<���<��<��<���<���<��<���<���<���<P��<���<���<���<9��<���<\��<��<I��<���<m��<޼�<`   `   ޼�<;��<��<d��<���<-��<���<���<d��<���<q��<��<��<{��<��<K��<���<���<F��<v��<U��<��<;��<μ�<`   `   ���<��<6��<-��<��<Y��<���<r��<��<��<���<��<���<��<��<r��<���<Y��<��<-��<)��<��<���<���<`   `   ���<d��<-��<��<N��<��<���<R��<=��<$��<���<���<��<%��<f��<���<���<+��<*��<J��<U��<���< ��< ��<`   `   ��<���<��<N��<���<Y��<*��< ��<���<���<���<���<��< ��<���<Y��<��<N��<���<���<5��<���<���<���<`   `   ��<-��<Y��<��<Y��<���<��<��<���<���<���<��<��<*��<���<6��<���<u��<F��< ��<���<���<���<���<`   `   ���<���<���<���<*��<��<���<���<1��<F��<S��<���<���<��<:��<���<���<���<���<���<���<z��<z��<���<`   `   ���<���<r��<R��< ��<��<���<��<C��<+��<���<���<��<���<f��<���<���<���<e��<���<'��<6��<���<L��<`   `   ��<d��<��<=��<���<���<1��<C��<4��<C��<��<���<��<=��<���<d��<0��<���<���<���<���<���<���<���<`   `   ���<���<��<$��<���<���<F��<+��<C��<h��<���<���<��<)��<��<���<M��<7��<#��<|��<m��<
��<8��<g��<`   `   ���<q��<���<���<���<���<S��<���<��<���<���<���<���<q��<���<>��<���<���<���<� �<���<���<p��<>��<`   `   ���<��<��<���<���<��<���<���<���<���<���<0��<��<y��<q��< �<��<��<m	�<T	�<��<�< �<^��<`   `   P��<��<���<��<��<��<���<��<��<��<���<��<f��<���<��<�	�<��<��<��<��<��<�	�<��<���<`   `   ���<{��<��<%��< ��<*��<��<���<=��<)��<q��<y��<���<�<?�<�<��<g�<��<��<��<+�<�<���<`   `   ���<��<��<f��<���<���<:��<f��<���<��<���<q��<��<?�<�<��<��<;�<��<��<0�<?�<��<q��<`   `   ���<K��<r��<���<Y��<6��<���<���<d��<���<>��< �<�	�<�<��<'�<� �<� �<@�<��<��<�	�< �<G��<`   `   9��<���<���<���<��<���<���<���<0��<M��<���<��<��<��<��<� �<�!�<� �<��<��<��<��<���<M��<`   `   ���<���<Y��<+��<N��<u��<���<���<���<7��<���<��<��<g�<;�<� �<� �<'�<��<�<��<��<8��<���<`   `   \��<F��<��<*��<���<F��<���<e��<���<#��<���<m	�<��<��<��<@�<��<��<w�<m	�<���<#��<���<e��<`   `   ��<v��<-��<J��<���< ��<���<���<���<|��<� �<T	�<��<��<��<��<��<�<m	�<� �<m��<���<���<���<`   `   I��<U��<)��<U��<5��<���<���<'��<���<m��<���<��<��<��<0�<��<��<��<���<m��<��<'��<h��<���<`   `   ���<��<��<���<���<���<z��<6��<���<
��<���<�<�	�<+�<?�<�	�<��<��<#��<���<'��<���<���<���<`   `   m��<;��<���< ��<���<���<z��<���<���<8��<p��< �<��<�<��< �<���<8��<���<���<h��<���<���< ��<`   `   ޼�<μ�<���< ��<���<���<���<L��<���<g��<>��<^��<���<���<q��<G��<M��<���<e��<���<���<���< ��<���<`   `   ?��<���<��<{��<���<���<���<���<��<}��<6��<)��<���<)��<��<}��<D��<���<g��<���<��<{��<���<���<`   `   ���<���<���<��<9��<���<���<���<Q��<���<<��<���<���<C��<���<;��<s��<���<���<��<��<���<���<���<`   `   ��<���<c��<O��<[��<���<p��<���<���<>��<(��<��<)��<>��<���<���<n��<���<a��<O��<[��<���<��<���<`   `   {��<��<O��<���<���<���<��<���<{��<U��<���<���<L��<e��<���<#��<���<���<��<i��<��<n��<���<���<`   `   ���<9��<[��<���<���<���<���<'��</��<���<��<���<N��<'��<���<���<���<���<&��<9��<���<^��<z��<^��<`   `   ���<���<���<���<���<���<��<���</��<���<���<��<���<+��<���<e��<���<���<���<���<���<I��<L��<���<`   `   ���<���<p��<��<���<��<���<��<���<4��<���<��<���<��<���<��<s��<���<���<���<{��<M��<g��<���<`   `   ���<���<���<���<'��<���<��<s��<:��<$��<l��<#��<���<��<���<���<s��<���<���<J��<T��<f��<M��<���<`   `   ��<Q��<���<{��</��</��<���<:��<`��<:��<���</��<Y��<{��<m��<Q��<;��<��<f��<���<���<���<~��<��<`   `   }��<���<>��<U��<���<���<4��<$��<:��<T��<���<���<L��<X��<���<p��<p��<���<���<���<���<s��<���<���<`   `   6��<<��<(��<���<��<���<���<l��<���<���<+��<���<��<<��<.��<���<���<��<i��<y��<���<��<���<���<`   `   )��<���<��<���<���<��<��<#��</��<���<���< ��<���<��<���<���<���<���<��<���<���<���<���<���<`   `   ���<���<)��<L��<N��<���<���<���<Y��<L��<��<���<	��<���<���<���<o �<��<��<��<e �<���<���<���<`   `   )��<C��<>��<e��<'��<+��<��<��<{��<X��<<��<��<���<���<��<��<��<��<�<��<��<���<���<���<`   `   ��<���<���<���<���<���<���<���<m��<���<.��<���<���<��<��<Z�<}�<�<E�<Z�<��<��<y��<���<`   `   }��<;��<���<#��<���<e��<��<���<Q��<p��<���<���<���<��<Z�<��<R�<o�< �<D�<��<���<���<���<`   `   D��<s��<n��<���<���<���<s��<s��<;��<p��<���<���<o �<��<}�<R�<��<R�<x�<��<x �<���<���<p��<`   `   ���<���<���<���<���<���<���<���<��<���<��<���<��<��<�<o�<R�<�<�<��<���<'��<���<���<`   `   g��<���<a��<��<&��<���<���<���<f��<���<i��<��<��<�<E�< �<x�<�<m�<��<t��<���<y��<���<`   `   ���<��<O��<i��<9��<���<���<J��<���<���<y��<���<��<��<Z�<D�<��<��<��<���<���<���<M��<���<`   `   ��<��<[��<��<���<���<{��<T��<���<���<���<���<e �<��<��<��<x �<���<t��<���< ��<T��<Y��<���<`   `   {��<���<���<n��<^��<I��<M��<f��<���<s��<��<���<���<���<��<���<���<'��<���<���<T��<l��<L��<=��<`   `   ���<���<��<���<z��<L��<g��<M��<~��<���<���<���<���<���<y��<���<���<���<y��<M��<Y��<L��<���<���<`   `   ���<���<���<���<^��<���<���<���<��<���<���<���<���<���<���<���<p��<���<���<���<���<=��<���<���<`   `   ,��<���<"��<���<���<���<3��<���<���<:��<���<���<W��<���<���<:��<���<���<���<���<)��<���<��<���<`   `   ���<���<<��<.��<���<���<���<s��<H��<���<���<���<���<���<���<6��<V��<��<���<���<��<R��<���<���<`   `   "��<<��<r��<:��<��<���<���<���<���<���<���<���<���<���<���<���<���<���<��<:��<n��<<��<'��<���<`   `   ���<.��<:��<���<c��<���<��<���<V��<���</��<3��<���<C��<���<4��<���<F��<���<P��<��<���<���<���<`   `   ���<���<��<c��<��<[��<c��<1��<��<p��<���<p��<$��<1��<0��<[��<H��<c��<���<���<��<���<���<���<`   `   ���<���<���<���<[��<:��<A��<���<���<S��<O��<���<���<]��<Q��<>��<���<���<���<z��<��<���<���</��<`   `   3��<���<���<��<c��<A��<���<U��<9��<���<P��<U��<���<A��<h��<��<���<���<!��<���<���<K��<u��<���<`   `   ���<s��<���<���<1��<���<U��<���<���<y��<���<q��<���<��<���<���<V��<���<_��<o��<9��<L��<t��<C��<`   `   ���<H��<���<V��<��<���<9��<���<���<���<"��<���</��<V��<���<H��<���<���<���<c��<���<c��<��<���<`   `   :��<���<���<���<p��<S��<���<y��<���<���<O��<T��<���<��<���<0��<
��<&��<���<��<��<���<+��<'��<`   `   ���<���<���</��<���<O��<P��<���<"��<O��<��</��<���<���<���<h��<���<��<`��<Z��<���<��<���<h��<`   `   ���<���<���<3��<p��<���<U��<q��<���<T��</��<���<���<���<���<���<��<7��<���<���<$��<-��<���<���<`   `   W��<���<���<���<$��<���<���<���</��<���<���<���<k��<���<���<���<���<���<x��<���<���<���<���<���<`   `   ���<���<���<C��<1��<]��<A��<��<V��<��<���<���<���<���<���<r��<o��<���<���<���<_��<���<���<���<`   `   ���<���<���<���<0��<Q��<h��<���<���<���<���<���<���<���<^��<��<I��<���<��<��<���<���<���<���<`   `   :��<6��<���<4��<[��<>��<��<���<H��<0��<h��<���<���<r��<��<���<_��<|��<���<��<_��<���<���<m��<`   `   ���<V��<���<���<H��<���<���<V��<���<
��<���<��<���<o��<I��<_��<M��<_��<E��<o��<���<��<���<
��<`   `   ���<��<���<F��<c��<���<���<���<���<&��<��<7��<���<���<���<|��<_��<���<���<���<$��< ��<+��<���<`   `   ���<���<��<���<���<���<!��<_��<���<���<`��<���<x��<���<��<���<E��<���<R��<���<n��<���<��<_��<`   `   ���<���<:��<P��<���<z��<���<o��<c��<��<Z��<���<���<���<��<��<o��<���<���<^��<��<P��<t��<��<`   `   )��<��<n��<��<��<��<���<9��<���<��<���<$��<���<_��<���<_��<���<$��<n��<��<���<9��<l��<��<`   `   ���<R��<<��<���<���<���<K��<L��<c��<���<��<-��<���<���<���<���<��< ��<���<P��<9��<g��<���<���<`   `   ��<���<'��<���<���<���<u��<t��<��<+��<���<���<���<���<���<���<���<+��<��<t��<l��<���<���<���<`   `   ���<���<���<���<���</��<���<C��<���<'��<h��<���<���<���<���<m��<
��<���<_��<��<��<���<���<���<`   `   ���<���<��<���<O��<Z��<o��<D��<&��<x��<���<���<*��<���<o��<x��<P��<D��<?��<Z��<y��<���<��<���<`   `   ���<\��<��<���<���<v��<k��<��<��<���<���<-��<"��<���<���<��<���<���<���<���<���<��<c��<���<`   `   ��<��<v��<K��<^��<��<���<?��<?��<Y��<���<a��<���<Y��<7��<?��<���<��<Z��<K��<x��<��<��<D��<`   `   ���<���<K��<-��<���<���<"��<���<��<���<���<���<���<	��<���<7��<���<���<H��<]��<���<���<���<���<`   `   O��<���<^��<���<_��<d��<���<e��<!��<���<���<���<:��<e��<\��<d��<���<���<2��<���<h��<���< ��<���<`   `   Z��<v��<��<���<d��<���<5��<���<7��<!��< ��<)��<���<K��<���<M��<���<���<���<S��<U��<���<���<h��<`   `   o��<k��<���<"��<���<5��<��<���<o��<G��<~��<���<��<5��<���<"��<���<k��<[��<���<��<W��<���<���<`   `   D��<��<?��<���<e��<���<���<:��<���<���<8��<���<���<N��<���<Q��<���<=��<���<���<	��<��<���<u��<`   `   &��<��<?��<��<!��<7��<o��<���<h��<���<[��<7��<C��<��<��<��<I��<���<���<��<���<��<���<���<`   `   x��<���<Y��<���<���<!��<G��<���<���<]��< ��<t��<���<j��<���<r��<U��<:��<��<}��<j��<���<A��<q��<`   `   ���<���<���<���<���< ��<~��<8��<[��< ��<���<���<���<���<x��<"��<Q��<���<W��<���<���<���<.��<"��<`   `   ���<-��<a��<���<���<)��<���<���<7��<t��<���<r��<"��<���<���<\��<o��<���<��< ��<���<���<c��<���<`   `   *��<"��<���<���<:��<���<��<���<C��<���<���<"��<<��<��<��<���<���<���<@��<���<���<���<��<��<`   `   ���<���<Y��<	��<e��<K��<5��<N��<��<j��<���<���<��<g��<v��<
��<���<w��<���<���<���<_��<n��<��<`   `   o��<���<7��<���<\��<���<���<���<��<���<w��<���<��<v��<O��<���<;��<"��<��<���<x��<v��<���<���<`   `   x��<��<?��<7��<d��<M��<"��<Q��<��<r��<"��<\��<���<
��<���<���<���<���<���<���<���<���<c��<#��<`   `   P��<���<���<���<���<���<���<���<I��<U��<Q��<o��<���<���<;��<���<��<���<7��<���<���<o��<I��<U��<`   `   D��<���<��<���<���<���<k��<=��<���<:��<���<���<���<w��<"��<���<���<��<���<���<���<���<A��<���<`   `   ?��<���<Z��<H��<2��<���<[��<���<���<��<W��<��<@��<���<��<���<7��<���<��<��<h��<��<���<���<`   `   Z��<���<K��<]��<���<S��<���<���<��<}��<���< ��<���<���<���<���<���<���<��<���<j��<��<���<���<`   `   y��<���<x��<���<h��<U��<��<	��<���<j��<���<���<���<���<x��<���<���<���<h��<j��<
��<	��<���<U��<`   `   ���<��<��<���<���<���<W��<��<��<���<���<���<���<_��<v��<���<o��<���<��<��<	��<m��<���<���<`   `   ��<c��<��<���< ��<���<���<���<���<A��<.��<c��<��<n��<���<c��<I��<A��<���<���<���<���<0��<���<`   `   ���<���<D��<���<���<h��<���<u��<���<q��<"��<���<��<��<���<#��<U��<���<���<���<U��<���<���<U��<`   `   ��<���<���<9��<��<��<+��<���<���<^��<b��<���<���<���<N��<^��<���<���<��<��<2��<9��<���<���<`   `   ���<���<���<���<o��<)��<V��<���<���<7��<f��<���<���<e��<K��<���<���<f��<A��<_��<���<���<���<���<`   `   ���<���< ��<���<���<���<?��<@��<e��<��<���<���<���<��<Z��<@��<I��<���<���<���<��<���<���<\��<`   `   9��<���<���<���<���<g��<���<T��<B��<;��<5��<5��</��<9��<i��<���<N��<���<���<���<���<6��<���<���<`   `   ��<o��<���<���<���<���<}��<���<���<���<���<���<���<���<Z��<���<���<���<o��<o��<$��<���<���<���<`   `   ��<)��<���<g��<���<��<���<���<��<_��<`��<���<���<���<!��<���<N��<��<A��<��< ��<���<���<��<`   `   +��<V��<?��<���<}��<���<���<Z��<���<���<���<Z��<���<���<y��<���<L��<V��<��<C��<(��<C��<��<C��<`   `   ���<���<@��<T��<���<���<Z��<T��<N��<E��<U��<j��<���<���<i��<K��<���<���<���<i��<j��<{��<q��<���<`   `   ���<���<e��<B��<���<��<���<N��<X��<N��<���<��<���<B��<E��<���<���<U��<��<<��<��<<��< ��<U��<`   `   ^��<7��<��<;��<���<_��<���<E��<N��<���<`��<���</��<)��<K��<[��<���<&��<|��<���<n��<d��<.��<���<`   `   b��<f��<���<5��<���<`��<���<U��<���<`��<���<5��<���<f��<P��<v��<���<o��<��<���<G��<o��<���<v��<`   `   ���<���<���<5��<���<���<Z��<j��<��<���<5��<��<���<���<���<;��<���<���<���<���<���<���<C��<���<`   `   ���<���<���</��<���<���<���<���<���</��<���<���<���<;��<r��<��<9��<l��<���<l��<1��<��<~��<;��<`   `   ���<e��<��<9��<���<���<���<���<B��<)��<f��<���<;��<���<���<���<��<B��<Z��<8��<���<���<���<G��<`   `   N��<K��<Z��<i��<Z��<!��<y��<i��<E��<K��<P��<���<r��<���<���<���<���<���<���<���<���<���<^��<���<`   `   ^��<���<@��<���<���<���<���<K��<���<[��<v��<;��<��<���<���<��<3��<K��<.��<q��<���<��<C��<u��<`   `   ���<���<I��<N��<���<N��<L��<���<���<���<���<���<9��<��<���<3��<��<3��<���<��<?��<���<���<���<`   `   ���<f��<���<���<���<��<V��<���<U��<&��<o��<���<l��<B��<���<K��<3��<���<Z��<x��<���<n��<.��<L��<`   `   ��<A��<���<���<o��<A��<��<���<��<|��<��<���<���<Z��<���<.��<���<Z��<v��<���<0��<|��<��<���<`   `   ��<_��<���<���<o��<��<C��<i��<<��<���<���<���<l��<8��<���<q��<��<x��<���<���<n��<3��<q��<R��<`   `   2��<���<��<���<$��< ��<(��<j��<��<n��<G��<���<1��<���<���<���<?��<���<0��<n��</��<j��<��< ��<`   `   9��<���<���<6��<���<���<C��<{��<<��<d��<o��<���<��<���<���<��<���<n��<|��<3��<j��<R��<���<���<`   `   ���<���<���<���<���<���<��<q��< ��<.��<���<C��<~��<���<^��<C��<���<.��<��<q��<��<���<���<���<`   `   ���<���<\��<���<���<��<C��<���<U��<���<v��<���<;��<G��<���<u��<���<L��<���<R��< ��<���<���<g��<`   `   ���<���<���<���<���<���<x��<���<��<���<���<��<���<��<���<���<7��<���<\��<���<���<���<���<���<`   `   ���<���<���<S��<T��<���<'��<h��<���<���<��<��<��<��<���<���<T��<0��<���<J��<D��<���<���<���<`   `   ���<���<���<���<���<���<���<��<H��<��<���<��<���<��<;��<��<���<���<���<���<���<���<���<e��<`   `   ���<S��<���<g��<y��<|��<J��<���<���<N��<H��<E��<C��<���<���<S��<h��<p��<z��<���<D��<���<U��<M��<`   `   ���<T��<���<y��<���<���<F��<���<��<"��<i��<"��<��<���<-��<���<��<y��<���<T��<���<s��<���<s��<`   `   ���<���<���<|��<���<���<��<���<v��<���<���<r��<x��<'��<���<���<h��<���<���<���<��<I��<Q��<,��<`   `   x��<'��<���<J��<F��<��<���<,��<(��<���<)��<,��<���<��<?��<J��<���<'��<d��< ��<��<e��<���< ��<`   `   ���<h��<��<���<���<���<,��<b��<���<���<e��<5��<x��<���<���<��<T��<���<���<���<4��<C��<���<���<`   `   ��<���<H��<���<��<v��<(��<���<���<���<��<v��<��<���<1��<���<3��<���<I��<W��<5��<W��<T��<���<`   `   ���<���<��<N��<"��<���<���<���<���<���<���<��<C��<��<���<���<b��<+��<���<���<���<���<3��<v��<`   `   ���<��<���<H��<i��<���<)��<e��<��<���<o��<H��<���<��<���<���<���<���<���<���<��<���<s��<���<`   `   ��<��<��<E��<"��<r��<,��<5��<v��<��<H��<��<��<��<���<���<��<��<��<���<��<��<���<���<`   `   ���<��<���<C��<��<x��<���<x��<��<C��<���<��<���<d��<���<��<���<���<F��<���<���<��<��<d��<`   `   ��<��<��<���<���<'��<��<���<���<��<��<��<d��<���<���<F��<���<S��<g��<���<7��<w��<���<n��<`   `   ���<���<;��<���<-��<���<?��<���<1��<���<���<���<���<���<���<���<���<%��<_��<���<���<���<���<���<`   `   ���<���<��<S��<���<���<J��<��<���<���<���<���<��<F��<���<q��<F��<Z��<���<���<7��<)��<���<���<`   `   7��<T��<���<h��<��<h��<���<T��<3��<b��<���<��<���<���<���<F��<���<F��<���<���<���<��<���<b��<`   `   ���<0��<���<p��<y��<���<'��<���<���<+��<���<��<���<S��<%��<Z��<F��<��<g��< ��<��<���<3��<���<`   `   \��<���<���<z��<���<���<d��<���<I��<���<���<��<F��<g��<_��<���<���<g��<(��<��<���<���<E��<���<`   `   ���<J��<���<���<T��<���< ��<���<W��<���<���<���<���<���<���<���<���< ��<��<���<���<S��<���<��<`   `   ���<D��<���<D��<���<��<��<4��<5��<���<��<��<���<7��<���<7��<���<��<���<���<H��<4��<��<��<`   `   ���<���<���<���<s��<I��<e��<C��<W��<���<���<��<��<w��<���<)��<��<���<���<S��<4��<n��<Q��<j��<`   `   ���<���<���<U��<���<Q��<���<���<T��<3��<s��<���<��<���<���<���<���<3��<E��<���<��<Q��<���<U��<`   `   ���<���<e��<M��<s��<,��< ��<���<���<v��<���<���<d��<n��<���<���<b��<���<���<��<��<j��<U��<k��<`   `   ���<��<���<#��<���<S��<���<���<��<��<���<X��<���<X��<���<��<��<���<���<S��<���<#��<���<��<`   `   ��<I��<���<���<C��<i��<���<���<���<b��<��<A��<8��<	��<n��<���<���<���<v��<A��<���<���<P��<!��<`   `   ���<���<u��<"��<���<���<���<���<C��<���<���<���<���<���<7��<���<���<���<���<"��<��<���<���<���<`   `   #��<���<"��<u��<h��<
��<���</��<���<���<��<��<���<���<;��<���<���<f��<���<"��<���<&��<��<	��<`   `   ���<C��<���<h��<���<��<���<.��<P��<���<��<���<X��<.��<���<��<���<h��<���<C��<���<���<5��<���<`   `   S��<i��<���<
��<��<���<���<%��<��<��<��<��<��<���<���<��<���<���<v��<U��<c��<'��<.��<n��<`   `   ���<���<���<���<���<���<v��<���<���<���<���<���<|��<���<���<���<���<���<���<���<���<Q��<���<���<`   `   ���<���<���</��<.��<%��<���<���<���<���<���<���<��<+��<;��<���<���<���<���<��<��<��<#��<���<`   `   ��<���<C��<���<P��<��<���<���<���<���<���<��<[��<���<7��<���<��<k��<���<���<���<���<���<k��<`   `   ��<b��<���<���<���<��<���<���<���<���<��<���<���<���<n��<��<���< ��<\��<���<���<O��<'��<���<`   `   ���<��<���<��<��<��<���<���<���<��<��<��<���<��<���<v��<��<���<���<��<���<���<��<v��<`   `   X��<A��<���<��<���<��<���<���<��<���<��<���<8��<Z��<��<2��<���<D��<���<���<9��<���<9��<��<`   `   ���<8��<���<���<X��<��<|��<��<[��<���<���<8��<���<���<���<��<9��<���<e��<���<6��<��<���<���<`   `   X��<	��<���<���<.��<���<���<+��<���<���<��<Z��<���<���<���<��<���<���<���<���<��<���<���<���<`   `   ���<n��<7��<;��<���<���<���<;��<7��<n��<���<��<���<���<��<"��<���<���<���<"��</��<���<���<��<`   `   ��<���<���<���<��<��<���<���<���<��<v��<2��<��<��<"��<���<���<���<���<��<��<
��<9��<r��<`   `   ��<���<���<���<���<���<���<���<��<���<��<���<9��<���<���<���<���<���<���<���<<��<���<��<���<`   `   ���<���<���<f��<h��<���<���<���<k��< ��<���<D��<���<���<���<���<���<���<���<���<9��<���<'��<k��<`   `   ���<v��<���<���<���<v��<���<���<���<\��<���<���<e��<���<���<���<���<���<P��<���<���<\��<���<���<`   `   S��<A��<"��<"��<C��<U��<���<��<���<���<��<���<���<���<"��<��<���<���<���<��<���<���<#��<���<`   `   ���<���<��<���<���<c��<���<��<���<���<���<9��<6��<��</��<��<<��<9��<���<���<���<��<���<c��<`   `   #��<���<���<&��<���<'��<Q��<��<���<O��<���<���<��<���<���<
��<���<���<\��<���<��<T��<.��<���<`   `   ���<P��<���<��<5��<.��<���<#��<���<'��<��<9��<���<���<���<9��<��<'��<���<#��<���<.��<1��<��<`   `   ��<!��<���<	��<���<n��<���<���<k��<���<v��<��<���<���<��<r��<���<k��<���<���<c��<���<��<���<`   `   H��<���<���<���<\��<��<���<���<���<B��<%��<���<6��<���<#��<B��<���<���<���<��<^��<���<���<���<`   `   ���<���<P��<���<���<G��<���<���<T��<���<���<���<���<���<���<X��<���<���<M��<���<���<L��<���<���<`   `   ���<P��<a��<
��<���<Y��<���<���<)��<���<	��<���<��<���<��<���<���<Y��<���<
��<k��<P��<���<���<`   `   ���<���<
��<j��<���<���<���<S��<���<<��<���<���<7��<���<Y��<���<���<���<p��<��<���<���<$��<��<`   `   \��<���<���<���<U��<���<���<��<f��<���<���<���<h��<��<���<���<X��<���<���<���<]��<Y��<��<Y��<`   `   ��<G��<Y��<���<���<(��<��</��<4��<��<��<8��<*��<��<-��<���<���<V��<M��<��<��<���<���<��<`   `   ���<���<���<���<���<��<��<���<��<���<��<���<��<��<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<S��<��</��<���<x��<���<���<|��<���<*��<��<Y��<���<���<���<.��<6��<i��<o��<;��<(��<`   `   ���<T��<)��<���<f��<4��<��<���<A��<���<��<4��<h��<���<'��<T��<���<��<O��<;��<R��<;��<P��<��<`   `   B��<���<���<<��<���<��<���<���<���<���<��<���<7��<���<���<F��<���<��<L��<���<���<F��<��<���<`   `   %��<���<	��<���<���<��<��<|��<��<��<~��<���<��<���<��<���<^��<���<��<-��<��<���<S��<���<`   `   ���<���<���<���<���<8��<���<���<4��<���<���<���<���<���<��<���<���<���<!��<��<���<���<���<��<`   `   6��<���<��<7��<h��<*��<��<*��<h��<7��<��<���<7��<a��<8��<���<���<���<���<���<���<���<8��<a��<`   `   ���<���<���<���<��<��<��<��<���<���<���<���<a��<���<���<��<��<���<���<��<	��<���<���<f��<`   `   #��<���<��<Y��<���<-��<���<Y��<'��<���<��<��<8��<���<��<��<���<E��<���<��<)��<���<-��<��<`   `   B��<X��<���<���<���<���<���<���<T��<F��<���<���<���<��<��<���<���<���<���<��<	��<���<���<���<`   `   ���<���<���<���<X��<���<���<���<���<���<^��<���<���<��<���<���<��<���<���<��<���<���<]��<���<`   `   ���<���<Y��<���<���<V��<���<���<��<��<���<���<���<���<E��<���<���<?��<���<���<���<���<��<!��<`   `   ���<M��<���<p��<���<M��<���<.��<O��<L��<��<!��<���<���<���<���<���<���<���<!��<��<L��<F��<.��<`   `   ��<���<
��<��<���<��<���<6��<;��<���<-��<��<���<��<��<��<��<���<!��<(��<���<?��<;��<���<`   `   ^��<���<k��<���<]��<��<���<i��<R��<���<��<���<���<	��<)��<	��<���<���<��<���<T��<i��<���<��<`   `   ���<L��<P��<���<Y��<���<���<o��<;��<F��<���<���<���<���<���<���<���<���<L��<?��<i��<���<���<\��<`   `   ���<���<���<$��<��<���<���<;��<P��<��<S��<���<8��<���<-��<���<]��<��<F��<;��<���<���<��<$��<`   `   ���<���<���<��<Y��<��<���<(��<��<���<���<��<a��<f��<��<���<���<!��<.��<���<��<\��<$��<���<`   `   ���<���<���<V��<���<���<���<��<���<n��<{��<���<���<���<���<n��<���<��<���<���<���<V��<��<���<`   `   ���<~��<3��<t��<��<���<R��<���<���<���<���<?��<=��<���<���<���<���<J��<���<��<t��<+��<���<���<`   `   ���<3��<��<���<:��<���<_��<���<J��<6��<n��<���<s��<6��<D��<���<e��<���<3��<���<���<3��<���<]��<`   `   V��<t��<���<Q��<~��<(��<U��<���<��<���<���<���<���<$��<���<M��<*��<���<O��<���<t��<[��<x��<v��<`   `   ���<��<:��<~��<���<���<<��<���<���<���<���<���<���<���<E��<���<���<~��<C��<��<���<���<���<���<`   `   ���<���<���<(��<���<���<Q��<?��<���<u��<y��<���<>��<I��<���<��<*��<���<���<���<t��<���<���<s��<`   `   ���<R��<_��<U��<<��<Q��<o��<i��<v��<C��<k��<i��<x��<Q��<4��<U��<d��<R��<���<��<@��<���<=��<��<`   `   ��<���<���<���<���<?��<i��<\��<^��<e��<`��<`��<>��<���<���<���<���<$��<"��<���<��<��<���<$��<`   `   ���<���<J��<��<���<���<v��<^��<@��<^��<z��<���<���<��<S��<���<���<���<��<��<���<��<���<���<`   `   n��<���<6��<���<���<u��<C��<e��<^��<:��<y��<��<���</��<���<s��<c��<���<(��<���<���<*��<���<a��<`   `   {��<���<n��<���<���<y��<k��<`��<z��<y��<���<���<w��<���<v��< ��<:��<���<���<���<���<���<9��< ��<`   `   ���<?��<���<���<���<���<i��<`��<���<��<���<���<=��<���<n��<���<>��<���<���<���<���<<��<���<o��<`   `   ���<=��<s��<���<���<>��<x��<>��<���<���<w��<=��<���<���<���<���<��<7��<e��<7��<��<���<���<���<`   `   ���<���<6��<$��<���<I��<Q��<���<��</��<���<���<���<0��<���<|��<���<��<��<���<|��<���<2��<���<`   `   ���<���<D��<���<E��<���<4��<���<S��<���<v��<n��<���<���<���<���<P��<���<T��<���<���<���<���<n��<`   `   n��<���<���<M��<���<��<U��<���<���<s��< ��<���<���<|��<���<f��<���<���<e��<���<|��<���<���<���<`   `   ���<���<e��<*��<���<*��<d��<���<���<c��<:��<>��<��<���<P��<���<��<���<Q��<���<��<>��<;��<c��<`   `   ��<J��<���<���<~��<���<R��<$��<���<���<���<���<7��<��<���<���<���<���<��<9��<���<���<���<���<`   `   ���<���<3��<O��<C��<���<���<"��<��<(��<���<���<e��<��<T��<e��<Q��<��<e��<���<���<(��<���<"��<`   `   ���<��<���<���<��<���<��<���<��<���<���<���<7��<���<���<���<���<9��<���<���<���<��<���<��<`   `   ���<t��<���<t��<���<t��<@��<��<���<���<���<���<��<|��<���<|��<��<���<���<���<���<��<F��<t��<`   `   V��<+��<3��<[��<���<���<���<��<��<*��<���<<��<���<���<���<���<>��<���<(��<��<��<���<���<���<`   `   ��<���<���<x��<���<���<=��<���<���<���<9��<���<���<2��<���<���<;��<���<���<���<F��<���<���<x��<`   `   ���<���<]��<v��<���<s��<��<$��<���<a��< ��<o��<���<���<n��<���<c��<���<"��<��<t��<���<x��<V��<`   `   k��<���<���<(��<���<��<h��<���<`��<���<���<V��<F��<V��<���<���<M��<���<~��<��<���<(��<���<���<`   `   ���<���<)��<V��<���<��<���<���<<��<���<��<��<��<��<���<E��<���<���<��<���<\��<��<���<���<`   `   ���<)��<c��<q��<���<��<���<y��<���<s��<���<���<���<s��<���<y��<���<��<���<q��<g��<)��<���<���<`   `   (��<V��<q��<���<���<6��<���<���<���<���<��<��<��<���<���<���<@��<���<���<g��<\��<-��<���<���<`   `   ���<���<���<���<���<N��<���<���<���<(��<(��<(��<���<���<���<N��<���<���<���<���<���<s��<'��<s��<`   `   ��<��<��<6��<N��<}��<���<L��<���<���<���<���<O��<���<u��<[��<@��<��<��<��<��<���<���<��<`   `   h��<���<���<���<���<���<���<l��<[��<��<N��<l��<���<���<���<���<���<���<l��<���<���<L��<���<���<`   `   ���<���<y��<���<���<L��<l��<���<k��<s��<���<`��<O��<���<���<n��<���<���<���<2��<���<���<1��<���<`   `   `��<<��<���<���<���<���<[��<k��<���<k��<d��<���<���<���<���<<��<Q��<{��<���<���<��<���<���<{��<`   `   ���<���<s��<���<(��<���<��<s��<k��<���<���<5��<��<h��<���<���<6��<u��<y��<���<���<���<u��<,��<`   `   ���<��<���<��<(��<���<N��<���<d��<���<��<��<���<��<���<W��<���<���<��<=��<���<���<���<W��<`   `   V��<��<���<��<(��<���<l��<`��<���<5��<��<���<��<[��<���<d��<}��<���< ��<*��<���<s��<d��<���<`   `   F��<��<���<��<���<O��<���<O��<���<��<���<��<>��<���<���<"��<f��<u��<���<u��<j��<"��<���<���<`   `   V��<��<s��<���<���<���<���<���<���<h��<��<[��<���<#��<���<���<���<���<���<���<���<���<"��<���<`   `   ���<���<���<���<���<u��<���<���<���<���<���<���<���<���<���<��<��<;��<,��<��<���<���<���<���<`   `   ���<E��<y��<���<N��<[��<���<n��<<��<���<W��<d��<"��<���<��<���<_��<U��<���<��<���<��<d��<S��<`   `   M��<���<���<@��<���<@��<���<���<Q��<6��<���<}��<f��<���<��<_��<l��<_��<��<���<c��<}��<���<6��<`   `   ���<���<��<���<���<��<���<���<{��<u��<���<���<u��<���<;��<U��<_��<B��<���<s��<���<���<u��<���<`   `   ~��<��<���<���<���<��<l��<���<���<y��<��< ��<���<���<,��<���<��<���<���< ��<
��<y��<���<���<`   `   ��<���<q��<g��<���<��<���<2��<���<���<=��<*��<u��<���<��<��<���<s��< ��<:��<���<���<1��<���<`   `   ���<\��<g��<\��<���<��<���<���<��<���<���<���<j��<���<���<���<c��<���<
��<���<���<���<���<��<`   `   (��<��<)��<-��<s��<���<L��<���<���<���<���<s��<"��<���<���<��<}��<���<y��<���<���<@��<���<���<`   `   ���<���<���<���<'��<���<���<1��<���<u��<���<d��<���<"��<���<d��<���<u��<���<1��<���<���<��<���<`   `   ���<���<���<���<s��<��<���<���<{��<,��<W��<���<���<���<���<S��<6��<���<���<���<��<���<���<���<`   `   ��<x��<p��<���<
��<0��<���<B��<���<���<���<2��<,��<2��<��<���<~��<B��<���<0��<���<���<���<x��<`   `   x��<���<J��<���<D��<���<���<!��<s��<���<���<���<���<���<���<}��<3��<���<���<U��<���<=��<���<}��<`   `   p��<J��<���<���<+��<g��<���<;��<4��<G��<z��<T��<v��<G��<8��<;��<���<g��<,��<���<���<J��<n��<4��<`   `   ���<���<���<��<z��</��<���<��</��<?��<E��<C��<F��<9��<��<���<A��<���<
��<���<���<���<���<���<`   `   
��<D��<+��<z��<���<���<���<���<��<���<���<���<���<���<���<���<���<z��<H��<D��<���<-��<=��<-��<`   `   0��<���<g��</��<���<���<r��<���<���<���<���<���<���<b��<���<���<A��<Z��<���<5��<���<P��<L��<���<`   `   ���<���<���<���<���<r��<���<���<��<9��<���<���<��<r��<��<���<���<���<���<���<���<���<���<���<`   `   B��<!��<;��<��<���<���<���<���<���<���<���<���<���<���<��</��<3��<G��<\��<[��<;��</��<X��<m��<`   `   ���<s��<4��</��<��<���<��<���<?��<���<��<���<���</��<O��<s��<���<���<j��<���<���<���<]��<���<`   `   ���<���<G��<?��<���<���<9��<���<���<)��<���<���<F��<:��<���<���<���<��<���<���<���<��<��<���<`   `   ���<���<z��<E��<���<���<���<���<��<���<���<E��<���<���<���<4��<���<���<���<���<���<���<���<4��<`   `   2��<���<T��<C��<���<���<���<���<���<���<E��<H��<���<7��<x��<~��<���<��<���<��< ��<���<z��<���<`   `   ,��<���<v��<F��<���<���<��<���<���<F��<���<���< ��<y��<���<���<^��<W��<���<W��<d��<���<���<y��<`   `   2��<���<G��<9��<���<b��<r��<���</��<:��<���<7��<y��<A��<s��<E��<���<���<���<���<P��<���<>��<r��<`   `   ��<���<8��<��<���<���<��<��<O��<���<���<x��<���<s��<i��<���<��<!��<$��<���<O��<s��<���<x��<`   `   ���<}��<;��<���<���<���<���</��<s��<���<4��<~��<���<E��<���<"��<��<��<��<���<P��<���<z��<2��<`   `   ~��<3��<���<A��<���<A��<���<3��<���<���<���<���<^��<���<��<��<���<��<��<���<Y��<���<���<���<`   `   B��<���<g��<���<z��<Z��<���<G��<���<��<���<��<W��<���<!��<��<��</��<���<Q��< ��<���<��<���<`   `   ���<���<,��<
��<H��<���<���<\��<j��<���<���<���<���<���<$��<��<��<���<���<���<���<���<d��<\��<`   `   0��<U��<���<���<D��<5��<���<[��<���<���<���<��<W��<���<���<���<���<Q��<���<���<���<���<X��<w��<`   `   ���<���<���<���<���<���<���<;��<���<���<���< ��<d��<P��<O��<P��<Y��< ��<���<���<���<;��<���<���<`   `   ���<=��<J��<���<-��<P��<���</��<���<��<���<���<���<���<s��<���<���<���<���<���<;��<���<L��<=��<`   `   ���<���<n��<���<=��<L��<���<X��<]��<��<���<z��<���<>��<���<z��<���<��<d��<X��<���<L��<0��<���<`   `   x��<}��<4��<���<-��<���<���<m��<���<���<4��<���<y��<r��<x��<2��<���<���<\��<w��<���<=��<���<(��<`   `   ���<���<��<3��<a��<���<���<8��<r��<���<���<��<���<��<��<���<P��<8��<��<���<?��<3��<,��<���<`   `   ���<��<���<J��<Z��<���<���<���<D��<���<���<���<���<���<���<O��<���<���<���<m��<Z��<���<���<���<`   `   ��<���<
��<���<4��<���<$��<)��<��<6��<���<s��<|��<6��<"��<)��<��<���<8��<���<��<���<��<���<`   `   3��<J��<���<z��<���<���<���<6��<��<2��<���<���<=��<"��<"��<���<���<���<c��<���<Z��<8��<��< ��<`   `   a��<Z��<4��<���<���<���<���<��< ��<#��<E��<#��<���<��<���<���<���<���<X��<Z��<L��<A��<���<A��<`   `   ���<���<���<���<���<;��<���<��<��<��<��<��<��<���<(��<
��<���<���<���<���<���<���<���<���<`   `   ���<���<$��<���<���<���<��<���<���<���<���<���<��<���<���<���<��<���<���<���< ��<��<��<���<`   `   8��<���<)��<6��<��<��<���<���<���<���<���<���<��<!��<"��<��<���<=��<M��<-��<7��<'��<'��<d��<`   `   r��<D��<��<��< ��<��<���<���<���<���<���<��<���<��<;��<D��<V��<���<q��<���<���<���<`��<���<`   `   ���<���<6��<2��<#��<��<���<���<���<���<��<5��<=��<)��<���<���<w��<���<M��<	��<��<d��<���<_��<`   `   ���<���<���<���<E��<��<���<���<���<��<2��<���<���<���<��<2��<-��<a��<���<o��<\��<a��<K��<2��<`   `   ��<���<s��<���<#��<��<���<���<��<5��<���<e��<���<��<"��<���<���<���<���<���<���<���<���<5��<`   `   ���<���<|��<=��<���<��<��<��<���<=��<���<���<}��<��<c��<���<N��<"��<&��<"��<U��<���<V��<��<`   `   ��<���<6��<"��<��<���<���<!��<��<)��<���<��<��<���<��<��<F��<���<���<.��<$��<��<���<���<`   `   ��<���<"��<"��<���<(��<���<"��<;��<���<��<"��<c��<��<&��<|��<9��<���<g��<|��<��<��<t��<"��<`   `   ���<O��<)��<���<���<
��<���<��<D��<���<2��<���<���<��<|��<���<���<���<{��<���<$��<���<���<1��<`   `   P��<���<��<���<���<���<��<���<V��<w��<-��<���<N��<F��<9��<���<���<���<<��<F��<G��<���<4��<w��<`   `   8��<���<���<���<���<���<���<=��<���<���<a��<���<"��<���<���<���<���<���<���<��<���<`��<���<���<`   `   ��<���<8��<c��<X��<���<���<M��<q��<M��<���<���<&��<���<g��<{��<<��<���<F��<���<s��<M��<l��<M��<`   `   ���<m��<���<���<Z��<���<���<-��<���<	��<o��<���<"��<.��<|��<���<F��<��<���<n��<��<���<'��<���<`   `   ?��<Z��<��<Z��<L��<���< ��<7��<���<��<\��<���<U��<$��<��<$��<G��<���<s��<��<���<7��<��<���<`   `   3��<���<���<8��<A��<���<��<'��<���<d��<a��<���<���<��<��<���<���<`��<M��<���<7��< ��<���<T��<`   `   ,��<���<��<��<���<���<��<'��<`��<���<K��<���<V��<���<t��<���<4��<���<l��<'��<��<���<���<��<`   `   ���<���<���< ��<A��<���<���<d��<���<_��<2��<5��<��<���<"��<1��<w��<���<M��<���<���<T��<��<���<`   `   ���<l��<���<ؾ�<׾�<��<��<���<��<ѿ�<x��<���<��<���<���<ѿ�<ۿ�<���<��<��<���<ؾ�<���<l��<`   `   l��<g��<Z��<U��<���<��<��<6��<���<��<���<���<���<���<Ϳ�<���<R��<
��<��<ƾ�<h��<K��<_��<p��<`   `   ���<Z��<���<���<���<)��<���<<��<B��<տ�<��<[��<׿�<տ�<M��<<��<���<)��<���<���<���<Z��<���<S��<`   `   ؾ�<U��<���<-��<��<��<6��<p��<t��<f��<+��<+��<r��<���<Y��<#��<
��<)��<��<���<h��<ݾ�<ľ�<̾�<`   `   ׾�<���<���<��<پ�<��<��<V��<*��<[��<]��<[��<��<V��</��<��<���<��<̾�<���<���<־�<���<־�<`   `   ��<��<)��<��<��<V��<1��<��<^��<p��<p��<i��<)��<��<?��<��<
��<��<��<#��<
��<
��<��<���<`   `   ��<��<���<6��<��<1��<M��<>��<S��<���<H��<>��<S��<1��<	��<6��<���<��< ��<��<?��<��<Z��<��<`   `   ���<6��<<��<p��<V��<��<>��<���<I��<T��<���<,��<)��<j��<Y��<-��<R��<���<Z��<p��<;��<'��<h��<u��<`   `   ��<���<B��<t��<*��<^��<S��<I��<F��<I��<f��<^��<
��<t��<g��<���<��<ݿ�<���<Ͽ�<���<Ͽ�<y��<ݿ�<`   `   ѿ�<��<տ�<f��<[��<p��<���<T��<I��<���<p��<o��<r��<ƿ�<Ϳ�<ֿ�<ٿ�<%��<��<���<���<-��<��<���<`   `   x��<���<��<+��<]��<p��<H��<���<f��<p��<I��<+��<��<���<���<߿�<.��<��<��<=��<ڿ�<��<S��<߿�<`   `   ���<���<[��<+��<[��<i��<>��<,��<^��<o��<+��<M��<���<���<%��<c��<6��<��<���<���<��<��<[��<<��<`   `   ��<���<׿�<r��<��<)��<S��<)��<
��<r��<��<���<��<C��<o��<x��<���<���<���<���<���<x��<a��<C��<`   `   ���<���<տ�<���<V��<��<1��<j��<t��<ƿ�<���<���<C��<���<U��<���<t��<���<���<X��<���<l��<{��<7��<`   `   ���<Ϳ�<M��<Y��</��<?��<	��<Y��<g��<Ϳ�<���<%��<o��<U��<���<'��<���<A��<���<'��<���<U��<���<%��<`   `   ѿ�<���<<��<#��<��<��<6��<-��<���<ֿ�<߿�<c��<x��<���<'��<~��<���<���<c��<>��<���<k��<[��<߿�<`   `   ۿ�<R��<���<
��<���<
��<���<R��<��<ٿ�<.��<6��<���<t��<���<���<���<���<���<t��<���<6��<6��<ٿ�<`   `   ���<
��<)��<)��<��<��<��<���<ݿ�<%��<��<��<���<���<A��<���<���<X��<���<���<��<��<��<��<`   `   ��<��<���<��<̾�<��< ��<Z��<���<��<��<���<���<���<���<c��<���<���<���<���<���<��<���<Z��<`   `   ��<ƾ�<���<���<���<#��<��<p��<Ͽ�<���<=��<���<���<X��<'��<>��<t��<���<���<>��<���<ڿ�<h��<
��<`   `   ���<h��<���<h��<���<
��<?��<;��<���<���<ڿ�<��<���<���<���<���<���<��<���<���<���<;��<Y��<
��<`   `   ؾ�<K��<Z��<ݾ�<־�<
��<��<'��<Ͽ�<-��<��<��<x��<l��<U��<k��<6��<��<��<ڿ�<;��<��<��<��<`   `   ���<_��<���<ľ�<���<��<Z��<h��<y��<��<S��<[��<a��<{��<���<[��<6��<��<���<h��<Y��<��<u��<ľ�<`   `   l��<p��<S��<̾�<־�<���<��<u��<ݿ�<���<߿�<<��<C��<7��<%��<߿�<ٿ�<��<Z��<
��<
��<��<ľ�<D��<`   `   ��<ݻ�<ܻ�<���<5��<<��<L��<���<���<Ӽ�<��<:��<��<:��<��<Ӽ�<���<���<|��<<��<��<���<���<ݻ�<`   `   ݻ�<!��<+��<��<���<���<d��<\��<Ǽ�<��<ڼ�<޼�<��<ۼ�<׼�<Ҽ�<{��<P��<}��<���<!��<��<��<��<`   `   ܻ�<+��<9��<"��<!��<
��<���<~��<n��<^��<��<��<޼�<^��<{��<~��<���<
��<)��<"��<3��<+��<��<���<`   `   ���<��<"��<y��<F��<��<T��<̼�<���<~��<���<���<���<���<���<A��<1��<Z��<\��<��<!��<��<���<��<`   `   5��<���<!��<F��<���<���<2��<���<���<���<_��<���<���<���<^��<���<���<F��<M��<���<��<��<9��<��<`   `   <��<���<
��<��<���<~��<V��<i��<v��<���<���<���<w��<C��<f��<μ�<1��<���<}��<@��<��<e��<\��<׻�<`   `   L��<d��<���<T��<2��<V��<˼�<6��<n��<���<d��<6��<м�<V��<6��<T��<���<d��<d��<Y��<���<S��<���<Y��<`   `   ���<\��<~��<̼�<���<i��<6��<=��<`��<l��<=��<"��<w��<���<���<o��<{��<���<ּ�<��<˼�<���<���<��<`   `   ���<Ǽ�<n��<���<���<v��<n��<`��<��<`��<���<v��<|��<���<���<Ǽ�<���<���<l��<ڼ�</��<ڼ�<X��<���<`   `   Ӽ�<��<^��<~��<���<���<���<l��<`��<y��<���<���<���<O��<׼�<׼�<���<��<���<��<��<��<��<���<`   `   ��<ڼ�<��<���<_��<���<d��<=��<���<���<L��<���<��<ڼ�<���<��<G��<x��<���<���<Y��<x��<n��<��<`   `   :��<޼�<��<���<���<���<6��<"��<v��<���<���<��<��<>��<���<"��<+��<���<u��<���<���<��<��<���<`   `   ��<��<޼�<���<���<w��<м�<w��<|��<���<��<��<���<,��<A��<6��<)��<˽�<��<˽�<2��<6��<2��<,��<`   `   :��<ۼ�<^��<���<���<C��<V��<���<���<O��<ڼ�<>��<,��<k��<Ľ�<���<ǽ�<$��<��<���<���<ݽ�<b��<��<`   `   ��<׼�<{��<���<^��<f��<6��<���<���<׼�<���<���<A��<Ľ�<��<���<���<J��<��<���<���<Ľ�<X��<���<`   `   Ӽ�<Ҽ�<~��<A��<���<μ�<T��<o��<Ǽ�<׼�<��<"��<6��<���<���<���<��<��<ݽ�<ǽ�<���<(��<��<��<`   `   ���<{��<���<1��<���<1��<���<{��<���<���<G��<+��<)��<ǽ�<���<��<s��<��<���<ǽ�<!��<+��<P��<���<`   `   ���<P��<
��<Z��<F��<���<d��<���<���<��<x��<���<˽�<$��<J��<��<��<c��<��<���<���<y��<��<���<`   `   |��<}��<)��<\��<M��<}��<d��<ּ�<l��<���<���<u��<��<��<��<ݽ�<���<��<D��<u��<u��<���<j��<ּ�<`   `   <��<���<"��<��<���<@��<Y��<��<ڼ�<��<���<���<˽�<���<���<ǽ�<ǽ�<���<u��<���<��<��<���<F��<`   `   ��<!��<3��<!��<��<��<���<˼�</��<��<Y��<���<2��<���<���<���<!��<���<u��<��<��<˼�<���<��<`   `   ���<��<+��<��<��<e��<S��<���<ڼ�<��<x��<��<6��<ݽ�<Ľ�<(��<+��<y��<���<��<˼�<@��<\��<4��<`   `   ���<��<��<���<9��<\��<���<���<X��<��<n��<��<2��<b��<X��<��<P��<��<j��<���<���<\��<-��<���<`   `   ݻ�<��<���<��<��<׻�<Y��<��<���<���<��<���<,��<��<���<��<���<���<ּ�<F��<��<4��<���<���<`   `   ��<b��<`��<K��<���<���<���<��<��<2��<ݹ�<G��<a��<G��<���<2��<���<��<ٹ�<���<���<K��<x��<b��<`   `   b��<N��<`��<O��<���<չ�<��<���<��<R��<��<���<��<��<9��<+��<���<ֹ�<���<���<d��<Q��<E��<f��<`   `   `��<`��<͹�<X��<L��<ƹ�<K��<Թ�<��<Թ�<��<ֹ�<���<Թ�<��<Թ�<@��<ƹ�<U��<X��<ǹ�<`��<e��<ֹ�<`   `   K��<O��<X��<ù�<ʹ�<���<���<��<��<߹�<��<��<��<���<���<���<���<޹�<���<I��<d��<O��<���<���<`   `   ���<���<L��<ʹ�<���<���<���<ɹ�<ٹ�<��<���<��<���<ɹ�<Ĺ�<���<���<ʹ�<x��<���<���<���<E��<���<`   `   ���<չ�<ƹ�<���<���<��<���<���<ܹ�<���<���<��<���<���<��<Ϲ�<���<���<���<���<ع�<ɹ�<���<ù�<`   `   ���<��<K��<���<���<���<M��<ݹ�<��<
��<׹�<ݹ�<S��<���<���<���<<��<��<¹�<���<Թ�<���<��<���<`   `   ��<���<Թ�<��<ɹ�<���<ݹ�<���<��<��<���<ʹ�<���<޹�<���<Ź�<���<��<%��<߹�<���<���<ֹ�<B��<`   `   ��<��<��<��<ٹ�<ܹ�<��<��<���<��<���<ܹ�<���<��<��<��<���<'��<��<��</��<��<ܹ�<'��<`   `   2��<R��<Թ�<߹�<��<���<
��<��<��<���<���<'��<��<Ź�<9��<6��<-��<O��<W��<��<��<t��<F��<��<`   `   ݹ�<��<��<��<���<���<׹�<���<���<���<���<��<��<��<��<?��<d��<+��<R��<7��<!��<+��<���<?��<`   `   G��<���<ֹ�<��<��<��<ݹ�<ʹ�<ܹ�<'��<��<ȹ�<��<K��<@��<���<G��<��<s��<���<0��<*��<���<X��<`   `   a��<��<���<��<���<���<S��<���<���<��<��<��<O��<��<F��<���<���<���<j��<���<���<���<7��<��<`   `   G��<��<Թ�<���<ɹ�<���<���<޹�<��<Ź�<��<K��<��<K��<���<O��<���<���<޺�<l��<d��<Һ�<B��<���<`   `   ���<9��<��<���<Ĺ�<��<���<���<��<9��<��<@��<F��<���<���<պ�<���<a��<���<պ�<_��<���<]��<@��<`   `   2��<+��<Թ�<���<���<Ϲ�<���<Ź�<��<6��<?��<���<���<O��<պ�</��<���<w��<��<��<d��<���<���<?��<`   `   ���<���<@��<���<���<���<<��<���<���<-��<d��<G��<���<���<���<���<���<���<���<���<���<G��<m��<-��<`   `   ��<ֹ�<ƹ�<޹�<ʹ�<���<��<��<'��<O��<+��<��<���<���<a��<w��<���<y��<޺�<y��<0��<,��<F��<3��<`   `   ٹ�<���<U��<���<x��<���<¹�<%��<��<W��<R��<s��<j��<޺�<���<��<���<޺�<���<s��<=��<W��<��<%��<`   `   ���<���<X��<I��<���<���<���<߹�<��<��<7��<���<���<l��<պ�<��<���<y��<s��<8��<��<��<ֹ�<���<`   `   ���<d��<ǹ�<d��<���<ع�<Թ�<���</��<��<!��<0��<���<d��<_��<d��<���<0��<=��<��<��<���<��<ع�<`   `   K��<Q��<`��<O��<���<ɹ�<���<���<��<t��<+��<*��<���<Һ�<���<���<G��<,��<W��<��<���<���<���<ƹ�<`   `   x��<E��<e��<���<E��<���<��<ֹ�<ܹ�<F��<���<���<7��<B��<]��<���<m��<F��<��<ֹ�<��<���<9��<���<`   `   b��<f��<ֹ�<���<���<ù�<���<B��<'��<��<?��<X��<��<���<@��<?��<-��<3��<%��<���<ع�<ƹ�<���<ǹ�<`   `   Ͷ�<��<ж�<��<��<��<���<"��<���<d��<��<y��<���<y��<��<d��<t��<"��<,��<��<��<��<��<��<`   `   ��<��<ݶ�<ζ�<��<F��<���<��<?��<o��<���<G��<S��<���<Y��<J��<��<��<,��<��<��<ζ�<��<��<`   `   ж�<ݶ�<M��<��<��<
��<���<���<��<��<���<-��<���<��<��<���<���<
��<��<��<H��<ݶ�<Զ�<ɶ�<`   `   ��<ζ�<��<m��<.��<��<#��<S��<V��<��<��<��<��<b��<=��<��<��<A��<S��<��<��<��<��<���<`   `   ��<��<��<.��<���<��<,��<H��<$��<N��</��<N��<��<H��<U��<��<϶�<.��<��<��<���<(��<���<(��<`   `   ��<F��<
��<��<��<~��<��<��<V��<4��<4��<a��<��<���<g��<*��<��<���<,��<��<��<���<��<���<`   `   ���<���<���<#��<,��<��<"��</��<%��<߶�<��</��<(��<��</��<#��<��<���<��<��<O��<U��<j��<��<`   `   "��<��<���<S��<H��<��</��<"��<��<��<"��<��<��<[��<=��<��<��<&��<?��<��<`��<M��<��<Y��<`   `   ���<?��<��<V��<$��<V��<%��<��<ܶ�<��<8��<V��<��<V��<&��<?��<{��<p��<A��<���<���<���</��<p��<`   `   d��<o��<��<��<N��<4��<߶�<��<��<Ͷ�<4��<a��<��<q��<Y��<h��<X��<_��<ڷ�<T��<g��<���<W��<=��<`   `   ��<���<���<��</��<4��<��<"��<8��<4��<��<��<���<���<��<x��<`��<y��<˷�<���<���<y��<���<x��<`   `   y��<G��<-��<��<N��<a��</��<��<V��<a��<��<��<S��<~��<���<Ʒ�<÷�<���<6��<P��<̷�<���<���<���<`   `   ���<S��<���<��<��<��<(��<��<��<��<���<S��<���<��<���<Է�<��<���<���<���<��<Է�<~��<��<`   `   y��<���<��<b��<H��<���<��<[��<V��<q��<���<~��<��<���<���<���<Ʒ�<��<��<���<���<ַ�<��<ط�<`   `   ��<Y��<��<=��<U��<g��</��<=��<&��<Y��<��<���<���<���<���<)��<��<"��<7��<)��<���<���<���<���<`   `   d��<J��<���<��<��<*��<#��<��<?��<h��<x��<Ʒ�<Է�<���<)��<D��<��<ɷ�<*��<@��<���<ȷ�<���<x��<`   `   t��<��<���<��<϶�<��<��<��<{��<X��<`��<÷�<��<Ʒ�<��<��<���<��<��<Ʒ�<
��<÷�<h��<X��<`   `   "��<��<
��<A��<.��<���<���<&��<p��<_��<y��<���<���<��<"��<ɷ�<��<8��<��<���<̷�<y��<W��<{��<`   `   ,��<,��<��<S��<��<,��<��<?��<A��<ڷ�<˷�<6��<���<��<7��<*��<��<��<۷�<6��<���<ڷ�<>��<?��<`   `   ��<��<��<��<��<��<��<��<���<T��<���<P��<���<���<)��<@��<Ʒ�<���<6��<���<g��<���<��<���<`   `   ��<��<H��<��<���<��<O��<`��<���<g��<���<̷�<��<���<���<���<
��<̷�<���<g��<���<`��<i��<��<`   `   ��<ζ�<ݶ�<��<(��<���<U��<M��<���<���<y��<���<Է�<ַ�<���<ȷ�<÷�<y��<ڷ�<���<`��<C��<��<<��<`   `   ��<��<Զ�<��<���<��<j��<��</��<W��<���<���<~��<��<���<���<h��<W��<>��<��<i��<��<���<��<`   `   ��<��<ɶ�<���<(��<���<��<Y��<p��<=��<x��<���<��<ط�<���<x��<X��<{��<?��<���<��<<��<��<���<`   `   P��<i��<R��<���<R��<���<���<���<Ӵ�<���<��<ɴ�<���<ɴ�<���<���<���<���<Ӵ�<���<1��<���<e��<i��<`   `   i��<���<]��<J��<���<���<t��<���<ݴ�<Ŵ�<���<���<���<���<���<��<Ǵ�<c��<޴�<Ѵ�<Z��<O��<���<n��<`   `   R��<]��<}��<W��<M��<A��<ڴ�<���<���<���<��<��<ش�<���<���<���<Դ�<A��<Q��<W��<{��<]��<S��<���<`   `   ���<J��<W��<o��<~��<{��<���<���<���<d��<���<���<m��<���<���<|��<���<���<Y��<I��<Z��<���<{��<���<`   `   R��<���<M��<~��<��<���<T��<Ҵ�<���<���<Ǵ�<���<���<Ҵ�<x��<���<���<~��<p��<���<>��<���<���<���<`   `   ���<���<A��<{��<���<���<���<���<���<���<���<���<���<���<w��<ɴ�<���<3��<޴�<���<(��<���<���<��<`   `   ���<t��<ڴ�<���<T��<���<��<z��<���<���<���<z��<��<���<U��<���<Ѵ�<t��<���<���<���<~��<մ�<���<`   `   ���<���<���<���<Ҵ�<���<z��<���<ش�<��<���<i��<���<��<���<���<Ǵ�<���<ߴ�<˴�<s��<c��<Ŵ�<���<`   `   Ӵ�<ݴ�<���<���<���<���<���<ش�<���<ش�<���<���<���<���<���<ݴ�<���<���<��<���<ʹ�<���<o��<���<`   `   ���<Ŵ�<���<d��<���<���<���<��<ش�<���<���<´�<m��<{��<���<ô�<���<ٴ�<ٴ�<���<Ŵ�<��<Ӵ�<���<`   `   ��<���<��<���<Ǵ�<���<���<���<���<���<���<���<��<���<���<&��<���<��<д�<���<���<��<��<&��<`   `   ɴ�<���<��<���<���<���<z��<i��<���<´�<���<��<���<δ�<&��<ƴ�<ش�<ܴ�<��< ��<��<���<���<8��<`   `   ���<���<ش�<m��<���<���<��<���<���<m��<��<���<y��<���<��<���<Y��<ϴ�<���<ϴ�<a��<���<s��<���<`   `   ɴ�<���<���<���<Ҵ�<���<���<��<���<{��<���<δ�<���<��</��<(��<��<2��<��<���<8��<A��<��<���<`   `   ���<���<���<���<x��<w��<U��<���<���<���<���<&��<��</��<8��<���<��<r��<��<���<��</��<���<&��<`   `   ���<��<���<|��<���<ɴ�<���<���<ݴ�<ô�<&��<ƴ�<���<(��<���<���<���<��<���<��<8��<���<���<%��<`   `   ���<Ǵ�<Դ�<���<���<���<Ѵ�<Ǵ�<���<���<���<ش�<Y��<��<��<���<���<���<��<��<S��<ش�<���<���<`   `   ���<c��<A��<���<~��<3��<t��<���<���<ٴ�<��<ܴ�<ϴ�<2��<r��<��<���<���<��<Ŵ�<��<��<Ӵ�<���<`   `   Ӵ�<޴�<Q��<Y��<p��<޴�<���<ߴ�<��<ٴ�<д�<��<���<��<��<���<��<��<���<��<���<ٴ�<z��<ߴ�<`   `   ���<Ѵ�<W��<I��<���<���<���<˴�<���<���<���< ��<ϴ�<���<���<��<��<Ŵ�<��<���<Ŵ�<���<Ŵ�<���<`   `   1��<Z��<{��<Z��<>��<(��<���<s��<ʹ�<Ŵ�<���<��<a��<8��<��<8��<S��<��<���<Ŵ�<���<s��<ִ�<(��<`   `   ���<O��<]��<���<���<���<~��<c��<���<��<��<���<���<A��</��<���<ش�<��<ٴ�<���<s��<m��<���<���<`   `   e��<���<S��<{��<���<���<մ�<Ŵ�<o��<Ӵ�<��<���<s��<��<���<���<���<Ӵ�<z��<Ŵ�<ִ�<���<���<{��<`   `   i��<n��<���<���<���<��<���<���<���<���<&��<8��<���<���<&��<%��<���<���<ߴ�<���<(��<���<{��<��<`   `   }��<���<���<��<#��<���<���<��<,��<	��<	��<Y��<���<Y��<��<	��<��<��<ұ�<���<��<��<��<���<`   `   ���<ձ�<б�<���<��<��<��<��<,��<g��<��<=��<D��<��<Y��<6��<��<��<��<��<��<ñ�<ұ�<��<`   `   ���<б�<F��<���<��<$��<L��<���<.��<7��<%��<��< ��<7��<1��<���<J��<$��<��<���<G��<б�<���<E��<`   `   ��<���<���<N��<=��<��<
��</��<6��<F��<��<��<L��<@��<!��<���<��<M��<>��<��<��<��<߱�<��<`   `   #��<��<��<=��<��<��<��< ��<��<7��<��<7��<��< ��<��<��<ı�<=��<��<��<��<��<ı�<��<`   `   ���<��<$��<��<��<;��<��<���<��<���<���<��<��<���<.��<%��<��<��<��<���<��<��<��<��<`   `   ���<��<L��<
��<��<��<Z��<��<#��<��<��<��<b��<��< ��<
��<H��<��<���<��<H��<��<V��<��<`   `   ��<��<���</��< ��<���<��<��<���<��<��<���<��<��<!��<��<��<$��<��<Q��<��<��<N��<#��<`   `   ,��<,��<.��<6��<��<��<#��<���<[��<���<0��<��<���<6��<G��<,��<��<^��<��<?��<|��<?��<��<^��<`   `   	��<g��<7��<F��<7��<���<��<��<���<��<���<F��<L��<+��<Y��<��<"��<���<<��<{��<���<L��<���<��<`   `   	��<��<%��<��<��<���<��<��<0��<���<۱�<��<*��<��<��<��<o��<^��<T��<���<8��<^��<���<��<`   `   Y��<=��<��<��<7��<��<��<���<��<F��<��<��<D��<^��<Z��<i��<A��<:��<���<���<E��<0��<e��<h��<`   `   ���<D��< ��<L��<��<��<b��<��<���<L��<*��<D��<���<c��<���<}��<���<���<���<���<���<}��<���<c��<`   `   Y��<��<7��<@��< ��<���<��<��<6��<+��<��<^��<c��<���<���<4��<g��<���<���<V��<?��<���<���<]��<`   `   ��<Y��<1��<!��<��<.��< ��<!��<G��<Y��<��<Z��<���<���<.��<���<���<X��<���<���<��<���<���<Z��<`   `   	��<6��<���<���<��<%��<
��<��<,��<��<��<i��<}��<4��<���<A��<���<���<0��<Ʋ�<?��<w��<e��<	��<`   `   ��<��<J��<��<ı�<��<H��<��<��<"��<o��<A��<���<g��<���<���<Ʋ�<���<���<g��<���<A��<u��<"��<`   `   ��<��<$��<M��<=��<��<��<$��<^��<���<^��<:��<���<���<X��<���<���<f��<���<���<E��<\��<���<h��<`   `   ұ�<��<��<>��<��<��<���<��<��<<��<T��<���<���<���<���<0��<���<���<Ͳ�<���<J��<<��<��<��<`   `   ���<��<���<��<��<���<��<Q��<?��<{��<���<���<���<V��<���<Ʋ�<g��<���<���<���<���<I��<N��<ܱ�<`   `   ��<��<G��<��<��<��<H��<��<|��<���<8��<E��<���<?��<��<?��<���<E��<J��<���<g��<��<Z��<��<`   `   ��<ñ�<б�<��<��<��<��<��<?��<L��<^��<0��<}��<���<���<w��<A��<\��<<��<I��<��<ڱ�<��<��<`   `   ��<ұ�<���<߱�<ı�<��<V��<N��<��<���<���<e��<���<���<���<e��<u��<���<��<N��<Z��<��<���<߱�<`   `   ���<��<E��<��<��<��<��<#��<^��<��<��<h��<c��<]��<Z��<	��<"��<h��<��<ܱ�<��<��<߱�<9��<`   `   ���<|��<���<���<���<��<���<��<ܯ�<��<���<���<��<���<ů�<��<ɯ�<��<ԯ�<��<���<���<���<|��<`   `   |��<e��<���<z��<v��<���<¯�<z��<���<��<Ư�<���<���<ï�<ۯ�<���<���<���<���<���<���<���<d��<���<`   `   ���<���<ԯ�<}��<^��<���<̯�<���<~��<���<��<���<��<���<}��<���<ί�<���<[��<}��<د�<���<���<���<`   `   ���<z��<}��<���<���<���<���<��<���<���<ͯ�<ʯ�<���<���<ܯ�<���<���<���<���<s��<���<���<���<���<`   `   ���<v��<^��<���<a��<���<į�<���<���<ͯ�<���<ͯ�<|��<���<ׯ�<���<J��<���<q��<v��<���<���<t��<���<`   `   ��<���<���<���<���<ϯ�<���<���<կ�<���<���<ޯ�<���<��<ǯ�<˯�<���<���<���<��<���<���<���<���<`   `   ���<¯�<̯�<���<į�<���<���<���<���<���<���<���<���<���<���<���<̯�<¯�<ï�<���<���<���<���<���<`   `   ��<z��<���<��<���<���<���<���<̯�<կ�<���<���<���<���<ܯ�<z��<���<��<���<���<Ư�<���<���<���<`   `   ܯ�<���<~��<���<���<կ�<���<̯�<��<̯�<ȯ�<կ�<x��<���<���<���<̯�<���<���<ů�<���<ů�<���<���<`   `   ��<��<���<���<ͯ�<���<���<կ�<̯�<���<���<ٯ�<���<���<ۯ�<��<���<���<���<s��<y��<ï�<���<���<`   `   ���<Ư�<��<ͯ�<���<���<���<���<ȯ�<���<���<ͯ�<��<Ư�<���<���<���<ѯ�<��<���<د�<ѯ�<į�<���<`   `   ���<���<���<ʯ�<ͯ�<ޯ�<���<���<կ�<ٯ�<ͯ�<���<���<���<���<��<¯�<��<���<���<��<���<��<���<`   `   ��<���<��<���<|��<���<���<���<x��<���<��<���<ٯ�<���<ݯ�< ��<��<ݯ�<���<ݯ�<��< ��<֯�<���<`   `   ���<ï�<���<���<���<��<���<���<���<���<Ư�<���<���<���<ï�<ܯ�<į�<���<��<���<��<˯�<���<���<`   `   ů�<ۯ�<}��<ܯ�<ׯ�<ǯ�<���<ܯ�<���<ۯ�<���<���<ݯ�<ï�<��<��<���<���<���<��<��<ï�<��<���<`   `   ��<���<���<���<���<˯�<���<z��<���<��<���<��< ��<ܯ�<��<��<ϯ�<ů�<֯�<���<��<���<��<���<`   `   ɯ�<���<ί�<���<J��<���<̯�<���<̯�<���<���<¯�<��<į�<���<ϯ�<��<ϯ�<���<į�<���<¯�<���<���<`   `   ��<���<���<���<���<���<¯�<��<���<���<ѯ�<��<ݯ�<���<���<ů�<ϯ�<���<��<گ�<��<ί�<���<���<`   `   ԯ�<���<[��<���<q��<���<ï�<���<���<���<��<���<���<��<���<֯�<���<��<���<���<��<���<���<���<`   `   ��<���<}��<s��<v��<��<���<���<ů�<s��<���<���<ݯ�<���<��<���<į�<گ�<���<���<y��<ͯ�<���<x��<`   `   ���<���<د�<���<���<���<���<Ư�<���<y��<د�<��<��<��<��<��<���<��<��<y��<���<Ư�<���<���<`   `   ���<���<���<���<���<���<���<���<ů�<ï�<ѯ�<���< ��<˯�<ï�<���<¯�<ί�<���<ͯ�<Ư�<���<���<���<`   `   ���<d��<���<���<t��<���<���<���<���<���<į�<��<֯�<���<��<��<���<���<���<���<���<���<h��<���<`   `   |��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<x��<���<���<���<���<`   `   ���<'��<B��<L��<���<P��<@��<A��<*��<E��<\��<n��<G��<n��<b��<E��< ��<A��<K��<P��<��<L��<H��<'��<`   `   '��<L��</��<��<f��<-��<���<P��<X��<��<W��<<��<;��<T��<��<_��<S��<���<*��<o��<��<(��<N��<,��<`   `   B��</��<��<O��<Q��</��<]��<���<a��<3��<z��<K��<��<3��<\��<���<c��</��<K��<O��<	��</��<;��<¬�<`   `   L��<��<O��<6��<<��<U��<���<\��<k��<4��<A��<=��<3��<q��<Z��<���<X��<E��<4��<H��<��<Q��<a��<_��<`   `   ���<f��<Q��<<��<���<S��<ެ�<w��<.��<��<=��<��<)��<w��<��<S��<���<<��<[��<f��<���<)��<z��<)��<`   `   P��<-��</��<U��<S��<��<A��<t��<E��<F��<J��<L��<s��<9��<��<\��<X��<'��<*��<U��<	��<X��<Z��<��<`   `   @��<���<]��<���<ެ�<A��<X��<1��<<��<���<1��<1��<a��<A��<׬�<���<b��<���<>��<=��<.��<Z��<-��<=��<`   `   A��<P��<���<\��<w��<t��<1��<3��<,��<3��<7��<)��<s��<���<Z��<���<S��<F��<f��<K��<M��<L��<M��<i��<`   `   *��<X��<a��<k��<.��<E��<<��<,��<L��<,��<@��<E��<'��<k��<j��<X��<"��<9��<k��<���<F��<���<g��<9��<`   `   E��<��<3��<4��<��<F��<���<3��<,��<���<J��<��<3��<,��<��<J��<Q��<]��<���<l��<m��<���<_��<N��<`   `   \��<W��<z��<A��<=��<J��<1��<7��<@��<J��<0��<A��<���<W��<Y��<��<���<p��<���<���<���<p��<���<��<`   `   n��<<��<K��<=��<��<L��<1��<)��<E��<��<A��<C��<;��<s��<���<`��<A��<p��<���<���<q��<?��<b��<���<`   `   G��<;��<��<3��<)��<s��<a��<s��<'��<3��<���<;��<C��<���<z��<2��<x��<���<Y��<���<z��<2��<v��<���<`   `   n��<T��<3��<q��<w��<9��<A��<���<k��<,��<W��<s��<���<���<|��<���<���<���<���<���<���<~��<���<���<`   `   b��<��<\��<Z��<��<��<׬�<Z��<j��<��<Y��<���<z��<|��<խ�<}��<}��<���<���<}��<ҭ�<|��<w��<���<`   `   E��<_��<���<���<S��<\��<���<���<X��<J��<��<`��<2��<���<}��<F��<���<���<D��<��<���<3��<b��<{��<`   `    ��<S��<c��<X��<���<X��<b��<S��<"��<Q��<���<A��<x��<���<}��<���<���<���<~��<���<v��<A��<���<Q��<`   `   A��<���</��<E��<<��<'��<���<F��<9��<]��<p��<p��<���<���<���<���<���< ��<���<���<q��<l��<_��<@��<`   `   K��<*��<K��<4��<[��<*��<>��<f��<k��<���<���<���<Y��<���<���<D��<~��<���<[��<���<���<���<c��<f��<`   `   P��<o��<O��<H��<f��<U��<=��<K��<���<l��<���<���<���<���<}��<��<���<���<���<���<m��<���<M��<5��<`   `   ��<��<	��<��<���<	��<.��<M��<F��<m��<���<q��<z��<���<ҭ�<���<v��<q��<���<m��<?��<M��<4��<	��<`   `   L��<(��</��<Q��<)��<X��<Z��<L��<���<���<p��<?��<2��<~��<|��<3��<A��<l��<���<���<M��<R��<Z��<2��<`   `   H��<N��<;��<a��<z��<Z��<-��<M��<g��<_��<���<b��<v��<���<w��<b��<���<_��<c��<M��<4��<Z��<o��<a��<`   `   '��<,��<¬�<_��<)��<��<=��<i��<9��<N��<��<���<���<���<���<{��<Q��<@��<f��<5��<	��<2��<a��<���<`   `   ���<ݪ�<���<��<��<ڪ�<��<��<��<��<	��<��<��<��<	��<��<��<��<��<ڪ�<��<��<���<ݪ�<`   `   ݪ�<��<˪�<��<��<��<���<��<���<��<��<��<��<��<��<��<
��<���<��<��<��<Ǫ�<��<��<`   `   ���<˪�<��<��<��<��<��<��<���<��<���<��<���<��<��<��<	��<��<��<��<��<˪�<���<ݪ�<`   `   ��<��<��<���<٪�<��<��<ɪ�<��<$��<���<���<��<
��<ͪ�<��<��<ݪ�<���<��<��<��<۪�<ת�<`   `   ��<��<��<٪�<���<��<��<��<��<��<*��<��<��<��<��<��<���<٪�<��<��<��<٪�<���<٪�<`   `   ڪ�<��<��<��<��<Q��<��<ת�<��<��<��<��<Ӫ�<��<U��<��<��<��<��<ު�<5��<ת�<۪�<9��<`   `   ��<���<��<��<��<��<˪�<��<&��<��<��<��<Ӫ�<��<��<��<	��<���<��<��<0��<��<(��<��<`   `   ��<��<��<ɪ�<��<ת�<��<;��<��<��<?��<��<Ӫ�<��<ͪ�<��<
��< ��<��<̪�<��<��<Ъ�<��<`   `   ��<���<���<��<��<��<&��<��<���<��<&��<��<��<��<���<���<��<$��<��<���<��<���<��<$��<`   `   ��<��<��<#��<��<��<��<��<��<��<��<��<��<��<��<���<��<��<Ϊ�< ��<���<ʪ�<��<��<`   `   	��<��<���<���<*��<��<��<?��<&��<��<!��<���<���<��<��<ɪ�<)��<��<���<���<���<��<!��<ɪ�<`   `   ��<��<��<���<��<��<��<��<��<��<���<��<��<��<��<��<J��<��<��<��<��<N��<	��<ު�<`   `   ��<��<���<��<��<Ӫ�<Ӫ�<Ӫ�<��<��<���<��<��<��<��<.��<#��<!��<6��<!��<#��<.��<��<��<`   `   ��<��<��<
��<��<��<��<��<��<��<��<��<��<��<���<���<��<Ȫ�<̪�<��<��<���<��<��<`   `   	��<��<��<ͪ�<��<U��<��<ͪ�<���<��<��<��<��<���<ʪ�<��<��<���<��<��<Ӫ�<���<��<��<`   `   ��<��<��<��<��<��<��<��<���<���<ɪ�<��<.��<���<��<���<���<��<���<��<��<2��<	��<Ū�<`   `   ��<
��<	��<��<���<��<	��<
��<��<��<)��<J��<#��<��<��<���<���<���<��<��<#��<J��<)��<��<`   `   ��<���<��<ݪ�<٪�<��<���< ��<$��<��<��<��<!��<Ȫ�<���<��<���<���<̪�<%��<��<ު�<��<(��<`   `   ��<��<��<���<��<��<��<��<��<Ϊ�<���<��<6��<̪�<��<���<��<̪�<-��<��<���<Ϊ�<ߪ�<��<`   `   ڪ�<��<��<��<��<ު�<��<̪�<���< ��<���<��<!��<��<��<��<��<%��<��<���<���<���<Ъ�<��<`   `   ��<��<��<��<��<5��<0��<��<��<���<���<��<#��<��<Ӫ�<��<#��<��<���<���<��<��<0��<5��<`   `   ��<Ǫ�<˪�<��<٪�<ת�<��<��<���<ʪ�<��<N��<.��<���<���<2��<J��<ު�<Ϊ�<���<��<��<۪�<ݪ�<`   `   ���<��<���<۪�<���<۪�<(��<Ъ�<��<��<!��<	��<��<��<��<	��<)��<��<ߪ�<Ъ�<0��<۪�<���<۪�<`   `   ݪ�<��<ݪ�<ת�<٪�<9��<��<��<$��<��<ɪ�<ު�<��<��<��<Ū�<��<(��<��<��<5��<ݪ�<۪�<٪�<`   `   Q��<ʨ�<���<���<���<���<��<���<���<���<��<˨�<ʨ�<˨�<��<���<���<���<ި�<���<���<���<���<ʨ�<`   `   ʨ�<���<���<˨�<{��<���<֨�<���<���<ۨ�<���<��<ި�<���<��<���<���<ר�<���<z��<è�<���<���<ͨ�<`   `   ���<���<ݨ�<���<���<���<���<���<���<���<}��<٨�<���<���<���<���<���<���<���<���<��<���<���<��<`   `   ���<˨�<���<���<��<���<��<���<���<Ũ�<���<���<���<���<Ȩ�<��<���< ��<���<���<è�<���<���<���<`   `   ���<{��<���<��<���<���<���<���<���<���<���<���<¨�<���<��<���<���<��<���<{��<���<ި�<��<ި�<`   `   ���<���<���<���<���<C��<���<��<���<s��<v��<���<ڨ�<���<L��<���<���<���<���<���<���<���<���<ƨ�<`   `   ��<֨�<���<��<���<���<ݨ�<ʨ�<���<���<���<ʨ�<��<���<��<��<���<֨�<ܨ�<���<���<���<���<���<`   `   ���<���<���<���<���<��<ʨ�<j��<���<���<n��<ʨ�<ڨ�<���<Ȩ�<���<���<���<���<���<Ш�<٨�<���<���<`   `   ���<���<���<���<���<���<���<���<Ҩ�<���<���<���<Ĩ�<���<���<���<���<���<��<��<���<��<��<���<`   `   ���<ۨ�<���<Ũ�<���<s��<���<���<���<���<v��<���<���<���<��< ��<̨�<���<���<��<��<��<���<֨�<`   `   ��<���<}��<���<���<v��<���<n��<���<v��<���<���<���<���<��<Ψ�<���<���<��<ب�<��<���<���<Ψ�<`   `   ˨�<��<٨�<���<���<���<ʨ�<ʨ�<���<���<���<٨�<ި�<ͨ�<��<���<٨�<��<���<���<��<��<���<��<`   `   ʨ�<ި�<���<���<¨�<ڨ�<��<ڨ�<Ĩ�<���<���<ި�<Ψ�<Ǩ�<��<ܨ�<���<���<���<���<���<ܨ�<��<Ǩ�<`   `   ˨�<���<���<���<���<���<���<���<���<���<���<ͨ�<Ǩ�<���<���<���<��<��<��<���<���<��<���<ͨ�<`   `   ��<��<���<Ȩ�<��<L��<��<Ȩ�<���<��<��<��<��<���<���<���<��< ��<��<���<
��<���<٨�<��<`   `   ���<���<���<��<���<���<��<���<���< ��<Ψ�<���<ܨ�<���<���<���<��<��<���<���<���<��<���<˨�<`   `   ���<���<���<���<���<���<���<���<���<̨�<���<٨�<���<��<��<��<!��<��<��<��<���<٨�<���<̨�<`   `   ���<ר�<���< ��<��<���<֨�<���<���<���<���<��<���<��< ��<��<��<���<��<Ũ�<��<��<���<���<`   `   ި�<���<���<���<���<���<ܨ�<���<��<���<��<���<���<��<��<���<��<��<��<���<��<���<��<���<`   `   ���<z��<���<���<{��<���<���<���<��<��<ب�<���<���<���<���<���<��<Ũ�<���<ը�<��<��<���<���<`   `   ���<è�<��<è�<���<���<���<Ш�<���<��<��<��<���<���<
��<���<���<��<��<��<���<Ш�<���<���<`   `   ���<���<���<���<ި�<���<���<٨�<��<��<���<��<ܨ�<��<���<��<٨�<��<���<��<Ш�<���<���<ܨ�<`   `   ���<���<���<���<��<���<���<���<��<���<���<���<��<���<٨�<���<���<���<��<���<���<���<��<���<`   `   ʨ�<ͨ�<��<���<ި�<ƨ�<���<���<���<֨�<Ψ�<��<Ǩ�<ͨ�<��<˨�<̨�<���<���<���<���<ܨ�<���<��<`   `   \��<���<t��<{��<���<���<���<a��<r��<R��<e��<���<a��<���<[��<R��<���<a��<���<���<���<{��<i��<���<`   `   ���<���<���<���<���<���<���<��<���<Y��<���<���<���<���<f��<���<֦�<���<���<���<���<���<���<���<`   `   t��<���<e��<���<���<A��<o��<���<���<ڦ�<���<���<���<ڦ�<���<���<y��<A��<���<���<l��<���<m��<d��<`   `   {��<���<���<���<o��<���<���<Q��<���<���<���<���<���<���<^��<���<���<h��<���<���<���<|��<]��<W��<`   `   ���<���<���<o��<���<���<���<���<s��<���<���<���<~��<���<���<���<Ц�<o��<���<���<���<���<���<���<`   `   ���<���<A��<���<���<o��<���<���<���<���<���<���<���<���<|��<���<���<F��<���<���<a��<s��<y��<l��<`   `   ���<���<o��<���<���<���<x��<���<���<ئ�<���<���<z��<���<���<���<z��<���<���<���<{��<¦�<i��<���<`   `   a��<��<���<Q��<���<���<���<r��<���<���<u��<���<���<���<^��<���<֦�<b��<���<���<���<���<���<���<`   `   r��<���<���<���<s��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<i��<C��<i��<���<���<`   `   R��<Y��<ڦ�<���<���<���<ئ�<���<���<ަ�<���<���<���<ަ�<f��<R��<���<k��<W��<}��<q��<I��<q��<̦�<`   `   e��<���<���<���<���<���<���<u��<���<���<���<���<���<���<X��<���<���<z��<���<u��<���<z��<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<Ħ�<���<{��<���<���<���<���<`   `   a��<���<���<���<~��<���<z��<���<���<���<���<���<i��<���<���<q��<a��<���<���<���<]��<q��<���<���<`   `   ���<���<ڦ�<���<���<���<���<���<���<ަ�<���<���<���<���<d��<���<���<l��<{��<Ŧ�<���<W��<���<Ȧ�<`   `   [��<f��<���<^��<���<|��<���<^��<���<f��<X��<���<���<d��<���<���<���<s��<���<���<æ�<d��<���<���<`   `   R��<���<���<���<���<���<���<���<���<R��<���<���<q��<���<���<7��<���<���<E��<���<���<y��<���<���<`   `   ���<֦�<y��<���<Ц�<���<z��<֦�<���<���<���<���<a��<���<���<���<s��<���<���<���<d��<���<���<���<`   `   a��<���<A��<h��<o��<F��<���<b��<���<k��<z��<Ħ�<���<l��<s��<���<���<f��<{��<���<���<x��<q��<���<`   `   ���<���<���<���<���<���<���<���<���<W��<���<���<���<{��<���<E��<���<{��<���<���<���<W��<���<���<`   `   ���<���<���<���<���<���<���<���<i��<}��<u��<{��<���<Ŧ�<���<���<���<���<���<r��<q��<f��<���<���<`   `   ���<���<l��<���<���<a��<{��<���<C��<q��<���<���<]��<���<æ�<���<d��<���<���<q��<Q��<���<o��<a��<`   `   {��<���<���<|��<���<s��<¦�<���<i��<I��<z��<���<q��<W��<d��<y��<���<x��<W��<f��<���<Ȧ�<y��<���<`   `   i��<���<m��<]��<���<y��<i��<���<���<q��<���<���<���<���<���<���<���<q��<���<���<o��<y��<���<]��<`   `   ���<���<d��<W��<���<l��<���<���<���<̦�<���<���<���<Ȧ�<���<���<���<���<���<���<a��<���<]��<i��<`   `   ���<d��<���<���<R��<Z��<c��<Y��<e��<r��<¤�<���<;��<���<���<r��<~��<Y��<F��<Z��<k��<���<z��<d��<`   `   d��<7��<{��<W��<F��<5��<t��<���<z��<W��<Ĥ�<��<v��<Ĥ�<g��<s��<���<��<G��<9��<I��<���<=��<b��<`   `   ���<{��< ��<w��<���<���<f��<]��<��<V��<D��<S��<N��<V��<v��<]��<m��<���<���<w��<��<{��<���<���<`   `   ���<W��<w��<K��<,��<���<:��<A��<w��<X��<a��<`��<O��<q��<Q��<F��<���< ��<]��<��<I��<���<���<z��<`   `   R��<F��<���<,��<U��<[��<���<���<v��<s��<���<s��<���<���<m��<[��<t��<,��<���<F��<a��<a��<]��<a��<`   `   Z��<5��<���<���<[��<r��<���<T��<d��<B��<B��<]��<K��<���<���<O��<���<���<G��<X��<���<`��<e��<���<`   `   c��<t��<f��<:��<���<���<��<���<i��<'��<o��<���<��<���<���<:��<p��<t��<S��<���<t��<���<a��<���<`   `   Y��<���<]��<A��<���<T��<���<���<]��<V��<���<���<K��<���<Q��<f��<���<V��<u��<H��<Y��<f��<M��<c��<`   `   e��<z��<��<w��<v��<d��<i��<]��<|��<]��<]��<d��<���<w��<g��<z��<z��<���<���<s��<���<s��<���<���<`   `   r��<W��<V��<X��<s��<B��<'��<V��<]��<2��<B��<g��<O��<_��<g��<o��<���<}��<z��<���<��<h��<���<���<`   `   ¤�<Ĥ�<D��<a��<���<B��<o��<���<]��<B��<���<a��<D��<Ĥ�<���<|��<���<c��<Z��<d��<y��<c��<t��<|��<`   `   ���<��<S��<`��<s��<]��<���<���<d��<g��<a��<\��<v��<���<?��<v��<���<���<���<w��<���<Ƥ�<|��<0��<`   `   ;��<v��<N��<O��<���<K��<��<K��<���<O��<D��<v��<F��<t��<���<Ĥ�<j��<���<��<���<d��<Ĥ�<���<t��<`   `   ���<Ĥ�<V��<q��<���<���<���<���<w��<_��<Ĥ�<���<t��<���<���<���<���<D��<V��<���<���<{��<���<}��<`   `   ���<g��<v��<Q��<m��<���<���<Q��<g��<g��<���<?��<���<���<L��<���<ۤ�<���<���<���<h��<���<{��<?��<`   `   r��<s��<]��<F��<[��<O��<:��<f��<z��<o��<|��<v��<Ĥ�<���<���<Ϥ�<ä�<դ�<��<u��<���<ͤ�<|��<{��<`   `   ~��<���<m��<���<t��<���<p��<���<z��<���<���<���<j��<���<ۤ�<ä�<#��<ä�<٤�<���<n��<���<���<���<`   `   Y��<��<���< ��<,��<���<t��<V��<���<}��<c��<���<���<D��<���<դ�<ä�<s��<V��<���<���<c��<���<��<`   `   F��<G��<���<]��<���<G��<S��<u��<���<z��<Z��<���<��<V��<���<��<٤�<V��<Ҥ�<���<h��<z��<���<u��<`   `   Z��<9��<w��<��<F��<X��<���<H��<s��<���<d��<w��<���<���<���<u��<���<���<���<c��<��<l��<M��<���<`   `   k��<I��<��<I��<a��<���<t��<Y��<���<��<y��<���<d��<���<h��<���<n��<���<h��<��<���<Y��<c��<���<`   `   ���<���<{��<���<a��<`��<���<f��<s��<h��<c��<Ƥ�<Ĥ�<{��<���<ͤ�<���<c��<z��<l��<Y��<���<e��<U��<`   `   z��<=��<���<���<]��<e��<a��<M��<���<���<t��<|��<���<���<{��<|��<���<���<���<M��<c��<e��<c��<���<`   `   d��<b��<���<z��<a��<���<���<c��<���<���<|��<0��<t��<}��<?��<{��<���<��<u��<���<���<U��<���<���<`   `   ���<S��<L��<I��<_��<f��<���<���<;��<���<���<d��<}��<d��<���<���<Z��<���<���<f��<~��<I��<:��<S��<`   `   S��<1��<���<���<U��<9��<o��<Q��<l��<:��<;��<y��<p��<<��<K��<a��<<��<��<L��<D��<���<���<6��<N��<`   `   L��<���<g��<���<���<���<��<x��<���<<��<f��<���<n��<<��<���<x��<��<���<���<���<h��<���<L��<o��<`   `   I��<���<���<M��<c��<���<���<���<f��<���<���<���<���<[��<���<���<���<R��<a��<���<���<D��<L��<G��<`   `   _��<U��<���<c��<N��<H��<���<<��<��<t��<]��<t��<���<<��<j��<H��<t��<c��<s��<U��<r��<M��<���<M��<`   `   f��<9��<���<���<H��<��<X��<���<t��<���<���<j��<{��<i��</��<7��<���<���<L��<a��<��<d��<i��<���<`   `   ���<o��<��<���<���<X��<w��<���<V��<���<b��<���<o��<X��<���<���<��<o��<���<q��<T��<g��<A��<q��<`   `   ���<Q��<x��<���<<��<���<���<5��<o��<d��<3��<���<{��<+��<���<���<<��<���<[��<T��<���<���<Y��<G��<`   `   ;��<l��<���<f��<��<t��<V��<o��<ˢ�<o��<G��<t��<���<f��<���<l��<U��<B��<���<K��<%��<K��<���<B��<`   `   ���<:��<<��<���<t��<���<���<d��<o��<���<���<c��<���<I��<K��<��<@��<`��<}��<L��<>��<i��<e��<U��<`   `   ���<;��<f��<���<]��<���<b��<3��<G��<���<o��<���<b��<;��<���<o��<B��<���<r��<A��<���<���<)��<o��<`   `   d��<y��<���<���<t��<j��<���<���<t��<c��<���<���<p��<_��<N��<U��<V��<z��<N��<:��<k��<k��<Z��<>��<`   `   }��<p��<n��<���<���<{��<o��<{��<���<���<b��<p��<���<���<s��<o��<��<p��<���<p��<��<o��<��<���<`   `   d��<<��<<��<[��<<��<i��<X��<+��<f��<I��<;��<_��<���<W��<h��<���<z��<V��<j��<���<z��<W��<\��<���<`   `   ���<K��<���<���<j��</��<���<���<���<K��<���<N��<s��<h��<���<H��<x��<s��<P��<H��<���<h��<e��<N��<`   `   ���<a��<x��<���<H��<7��<���<���<l��<��<o��<U��<o��<���<H��<��<[��<p��<���<7��<z��<w��<Z��<p��<`   `   Z��<<��<��<���<t��<���<��<<��<U��<@��<B��<V��<��<z��<x��<[��<��<[��<u��<z��<��<V��<<��<@��<`   `   ���<��<���<R��<c��<���<o��<���<B��<`��<���<z��<p��<V��<s��<p��<[��<c��<j��<x��<k��<���<e��<7��<`   `   ���<L��<���<a��<s��<L��<���<[��<���<}��<r��<N��<���<j��<P��<���<u��<j��<z��<N��<~��<}��<���<[��<`   `   f��<D��<���<���<U��<a��<q��<T��<K��<L��<A��<:��<p��<���<H��<7��<z��<x��<N��<B��<>��<A��<Y��<���<`   `   ~��<���<h��<���<r��<��<T��<���<%��<>��<���<k��<��<z��<���<z��<��<k��<~��<>��<=��<���<?��<��<`   `   I��<���<���<D��<M��<d��<g��<���<K��<i��<���<k��<o��<W��<h��<w��<V��<���<}��<A��<���<w��<i��<;��<`   `   :��<6��<L��<L��<���<i��<A��<Y��<���<e��<)��<Z��<��<\��<e��<Z��<<��<e��<���<Y��<?��<i��<���<L��<`   `   S��<N��<o��<G��<M��<���<q��<G��<B��<U��<o��<>��<���<���<N��<p��<@��<7��<[��<���<��<;��<L��<|��<`   `   V��<t��<���<L��<���<}��<���<���<u��<q��<���<O��<|��<O��<l��<q��<���<���<Z��<}��<���<L��<t��<t��<`   `   t��<���<n��<���<y��<J��<���<���<g��<W��<u��<t��<m��<y��<h��<Y��<���<���<_��<d��<y��<��<���<m��<`   `   ���<n��<���<Q��<t��<a��<��<���<���<���<��<Z��<���<���<���<���<��<a��<u��<Q��<���<n��<���<���<`   `   L��<���<Q��<7��<q��<���<���<��<=��<���<<��<@��<���</��</��<���<q��<\��<K��<b��<y��<E��<g��<d��<`   `   ���<y��<t��<q��<_��<n��<���<(��<u��<*��<]��<*��<���<(��<p��<n��<���<q��<O��<y��<���<W��<Ǡ�<W��<`   `   }��<J��<a��<���<n��<���<���<���<D��<���<���<6��<���<���<���<Y��<q��<q��<_��<u��<l��<f��<j��<z��<`   `   ���<���<��<���<���<���<@��<g��<U��<���<f��<g��<3��<���<���<���<��<���<v��<P��<S��<P��<B��<P��<`   `   ���<���<���<��<(��<���<g��<l��<Y��<K��<h��<{��<���<��</��<���<���<���<0��<���<���<ɠ�<���<��<`   `   u��<g��<���<=��<u��<D��<U��<Y��<_��<Y��<D��<D��<���<=��<j��<g��<���<v��<���<|��<T��<|��<���<v��<`   `   q��<W��<���<���<*��<���<���<K��<Y��<Ġ�<���<��<���<Ϡ�<h��<i��<���<���<6��<���<{��<"��<���<���<`   `   ���<u��<��<<��<]��<���<f��<h��<D��<���<v��<<��<v��<u��<w��<���<���<v��<���<��<���<v��<i��<���<`   `   O��<t��<Z��<@��<*��<6��<g��<{��<D��<��<<��<k��<m��<H��<|��<���<���<���<l��<X��<���<���<���<l��<`   `   |��<m��<���<���<���<���<3��<���<���<���<v��<m��<���<���<���<���<a��<���<l��<���<Y��<���<���<���<`   `   O��<y��<���</��<(��<���<���<��<=��<Ϡ�<u��<H��<���<A��<G��<���<���<V��<k��<Ԡ�<���<6��<E��<���<`   `   l��<h��<���</��<p��<���<���</��<j��<h��<w��<|��<���<G��<���<���<���<q��<���<���<Ơ�<G��<���<|��<`   `   q��<Y��<���<���<n��<Y��<���<���<g��<i��<���<���<���<���<���<e��<���<Ԡ�<y��<���<���<���<���<���<`   `   ���<���<��<q��<���<q��<��<���<���<���<���<���<a��<���<���<���<���<���<���<���<g��<���<{��<���<`   `   ���<���<a��<\��<q��<q��<���<���<v��<���<v��<���<���<V��<q��<Ԡ�<���<`��<k��<���<���<z��<���<h��<`   `   Z��<_��<u��<K��<O��<_��<v��<0��<���<6��<���<l��<l��<k��<���<y��<���<k��<P��<l��<���<6��<���<0��<`   `   }��<d��<Q��<b��<y��<u��<P��<���<|��<���<��<X��<���<Ԡ�<���<���<���<���<l��<��<{��<o��<���<d��<`   `   ���<y��<���<y��<���<l��<S��<���<T��<{��<���<���<Y��<���<Ơ�<���<g��<���<���<{��<o��<���<<��<l��<`   `   L��<��<n��<E��<W��<f��<P��<ɠ�<|��<"��<v��<���<���<6��<G��<���<���<z��<6��<o��<���<d��<j��<B��<`   `   t��<���<���<g��<Ǡ�<j��<B��<���<���<���<i��<���<���<E��<���<���<{��<���<���<���<<��<j��<٠�<g��<`   `   t��<m��<���<d��<W��<z��<P��<��<v��<���<���<l��<���<���<|��<���<���<h��<0��<d��<l��<B��<g��<���<`   `   ���<n��<���<���<x��<���<���<N��<]��<{��<ў�<���<���<���<���<{��<���<N��<o��<���<���<���<}��<n��<`   `   n��<l��<���<���<b��<b��<���<���<`��<t��<���<���<���<���<���<P��<���<���<u��<J��<���<���<n��<d��<`   `   ���<���<l��<֞�<Ğ�<���<e��<���<���<���<K��<���<L��<���<���<���<c��<���<Ȟ�<֞�<f��<���<���<y��<`   `   ���<���<֞�<���<���<���<���<o��<���<o��<���<ƞ�<i��<���<��<���<���<w��<���<��<���<���<���<���<`   `   x��<b��<Ğ�<���<���<Z��<���<˞�<��<���<"��<���<���<˞�<x��<Z��<���<���<���<b��<���<d��<���<d��<`   `   ���<b��<���<���<Z��<e��<���<ʞ�<���<���<���<t��<Ğ�<���<u��<B��<���<Ϟ�<u��<{��<���<���<���<���<`   `   ���<���<e��<���<���<���<��<���<}��<?��<���<���<ߝ�<���<���<���<g��<���<���<̞�<���<���<x��<̞�<`   `   N��<���<���<o��<˞�<ʞ�<���<��<���<���<��<Ğ�<Ğ�<���<��<˞�<���<D��<m��<���<L��<Y��<���<Y��<`   `   ]��<`��<���<���<��<���<}��<���<ƞ�<���<l��<���<��<���<z��<`��<|��<~��<���<t��<s��<t��<͞�<~��<`   `   {��<t��<���<o��<���<���<?��<���<���<V��<���<n��<i��<���<���<q��<���<���<e��<ޞ�<ў�<Q��<���<���<`   `   ў�<���<K��<���<"��<���<���<��<l��<���<@��<���<>��<���<ʞ�<g��<Z��<���<O��<���<o��<���<D��<g��<`   `   ���<���<���<ƞ�<���<t��<���<Ğ�<���<n��<���<���<���<���<i��<S��<���<���<S��<?��<���<���<U��<Y��<`   `   ���<���<L��<i��<���<Ğ�<ߝ�<Ğ�<��<i��<>��<���<���<}��<���<���<V��<���<��<���<N��<���<���<}��<`   `   ���<���<���<���<˞�<���<���<���<���<���<���<���<}��<���<���<r��<i��<u��<���<~��<f��<���<���<���<`   `   ���<���<���<��<x��<u��<���<��<z��<���<ʞ�<i��<���<���<x��<N��<���<m��<x��<N��<���<���<���<i��<`   `   {��<P��<���<���<Z��<B��<���<˞�<`��<q��<g��<S��<���<r��<N��<���<���<���<���<?��<f��<���<U��<l��<`   `   ���<���<c��<���<���<���<g��<���<|��<���<Z��<���<V��<i��<���<���<���<���<���<i��<]��<���<S��<���<`   `   N��<���<���<w��<���<Ϟ�<���<D��<~��<���<���<���<���<u��<m��<���<���<]��<���<���<���<���<���<n��<`   `   o��<u��<Ȟ�<���<���<u��<���<m��<���<e��<O��<S��<��<���<x��<���<���<���<ў�<S��<V��<e��<ʞ�<m��<`   `   ���<J��<֞�<��<b��<{��<̞�<���<t��<ޞ�<���<?��<���<~��<N��<?��<i��<���<S��<���<ў�<d��<���<��<`   `   ���<���<f��<���<���<���<���<L��<s��<ў�<o��<���<N��<f��<���<f��<]��<���<V��<ў�<���<L��<n��<���<`   `   ���<���<���<���<d��<���<���<Y��<t��<Q��<���<���<���<���<���<���<���<���<e��<d��<L��<���<���<L��<`   `   }��<n��<���<���<���<���<x��<���<͞�<���<D��<U��<���<���<���<U��<S��<���<ʞ�<���<n��<���<���<���<`   `   n��<d��<y��<���<d��<���<̞�<Y��<~��<���<g��<Y��<}��<���<i��<l��<���<n��<m��<��<���<L��<���<���<`   `   ?��<�<���<Μ�<���<���<���<ڜ�<��<ל�<��<���<���<���<Ԝ�<ל�<��<ڜ�<Ӝ�<���<ڜ�<Μ�<���<�<`   `   �<���<Ɯ�<���<���<���<���<��<���<���<���<Ĝ�<���<���<���<���<М�<Ϝ�<���<r��<���<ڜ�<���<���<`   `   ���<Ɯ�<���<���<ݜ�<˜�<E��<؜�<��<М�<���<��<���<М�<��<؜�<@��<˜�<��<���<y��<Ɯ�<���<���<`   `   Μ�<���<���<F��<s��<ޜ�<Ϝ�<���<���<Ɯ�<���<Ŝ�<���<���<���<��<̜�<Z��<X��<Μ�<���<Ü�<Ҝ�<ќ�<`   `   ���<���<ݜ�<s��<��<̜�<ќ�<o��<���<s��<|��<s��<���<o��<���<̜�<��<s��<���<���<̜�<���<���<���<`   `   ���<���<˜�<ޜ�<̜�<���<��<���<���<Ԝ�<Μ�<���<���<���<���<���<̜�<ߜ�<���<���<���<���<���<���<`   `   ���<���<E��<Ϝ�<ќ�<��<���<Ȝ�<���<
��<˜�<Ȝ�<���<��<ܜ�<Ϝ�<D��<���<���<Ԝ�<���<)��<~��<Ԝ�<`   `   ڜ�<��<؜�<���<o��<���<Ȝ�<f��<���<���<`��<���<���<V��<���<��<М�<Ϝ�<ڜ�<���<��<���<���<Ȝ�<`   `   ��<���<��<���<���<���<���<���<��<���<���<���<���<���<Ü�<���<���<���<Ӝ�<���<ɜ�<���<��<���<`   `   ל�<���<М�<Ɯ�<s��<Ԝ�<
��<���<���<"��<Μ�<Y��<���<��<���<̜�<͜�<���<Ӝ�<���<���<���<���<ߜ�<`   `   ��<���<���<���<|��<Μ�<˜�<`��<���<Μ�<���<���<���<���<��<��<���<��<ʜ�<���<��<��<���<��<`   `   ���<Ĝ�<��<Ŝ�<s��<���<Ȝ�<���<���<Y��<���<��<���<���<М�<̜�<���<��<М�<���<ڜ�<��<͜�<�<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<Ü�<���<Ɯ�<���<���<��<���<���<Ɯ�<ʜ�<Ü�<`   `   ���<���<М�<���<o��<���<��<V��<���<��<���<���<Ü�<���<���<��<��<���<���<��<��<���<���<Ȝ�<`   `   Ԝ�<���<��<���<���<���<ܜ�<���<Ü�<���<��<М�<���<���<��<ۜ�<���<՜�<Ϝ�<ۜ�<��<���<���<М�<`   `   ל�<���<؜�<��<̜�<���<Ϝ�<��<���<̜�<��<̜�<Ɯ�<��<ۜ�<���<��<��<���<͜�<��<ʜ�<͜�<��<`   `   ��<М�<@��<̜�<��<̜�<D��<М�<���<͜�<���<���<���<��<���<��<���<��<��<��<���<���<���<͜�<`   `   ڜ�<Ϝ�<˜�<Z��<s��<ߜ�<���<Ϝ�<���<���<��<��<���<���<՜�<��<��<ǜ�<���<���<ڜ�<��<���<���<`   `   Ӝ�<���<��<X��<���<���<���<ڜ�<Ӝ�<Ӝ�<ʜ�<М�<��<���<Ϝ�<���<��<���<���<М�<Ϝ�<Ӝ�<��<ڜ�<`   `   ���<r��<���<Μ�<���<���<Ԝ�<���<���<���<���<���<���<��<ۜ�<͜�<��<���<М�<���<���<���<���<��<`   `   ڜ�<���<y��<���<̜�<���<���<��<ɜ�<���<��<ڜ�<���<��<��<��<���<ڜ�<Ϝ�<���<��<��<q��<���<`   `   Μ�<ڜ�<Ɯ�<Ü�<���<���<)��<���<���<���<��<��<Ɯ�<���<���<ʜ�<���<��<Ӝ�<���<��<A��<���<���<`   `   ���<���<���<Ҝ�<���<���<~��<���<��<���<���<͜�<ʜ�<���<���<͜�<���<���<��<���<q��<���<ǜ�<Ҝ�<`   `   �<���<���<ќ�<���<���<Ԝ�<Ȝ�<���<ߜ�<��<�<Ü�<Ȝ�<М�<��<͜�<���<ڜ�<��<���<���<Ҝ�<Μ�<`   `   ���<ۚ�<ݚ�<���<:��<��<Ӛ�<ۚ�<��<˚�<��<��<���<��<ߚ�<˚�<��<ۚ�<���<��<[��<���<ɚ�<ۚ�<`   `   ۚ�<0��<��<��< ��<К�<��<-��<њ�<��<��<��<��<"��<���<���<��<+��<���<��<���<,��<0��<К�<`   `   ݚ�<��<ʚ�<��<W��<%��<���<���<���<1��<��<���<ߚ�<1��<���<���<���<%��<`��<��<���<��<��<��<`   `   ���<��<��<
��<��<��<��<��<��<V��<���<��<S��<ޚ�<���<1��<���<��<��<(��<���<���<���<���<`   `   :��< ��<W��<��<��<Ě�<'��<֚�</��<$��<���<$��<D��<֚�<��<Ě�<:��<��<3��< ��<N��< ��<"��< ��<`   `   ��<К�<%��<��<Ě�<���<)��<��<��<��<��<��<��<@��<���<���<���<9��<���<ޚ�<$��<��<��<-��<`   `   Ӛ�<��<���<��<'��<)��<��<&��<���</��<��<&��<��<)��<4��<��<���<��<Ϛ�<���<���<���<���<���<`   `   ۚ�<-��<���<��<֚�<��<&��<Ӛ�<��<ښ�<˚�<=��<��<���<���<��<��<К�<��<���<��<��<���<ݚ�<`   `   ��<њ�<���<��</��<��<���<��<{��<��<��<��<K��<��<ؚ�<њ�<��<ך�<,��<��<��<��<<��<ך�<`   `   ˚�<��<1��<V��<$��<��</��<ښ�<��<F��<��<��<S��<E��<���<���<��<Ț�<��<���<��<ݚ�<Ț�<��<`   `   ��<��<��<���<���<��<��<˚�<��<��<֚�<���<Қ�<��<��<��<ޚ�<Ϛ�<��<��<��<Ϛ�<Κ�<��<`   `   ��<��<���<��<$��<��<&��<=��<��<��<���<��<��<��<��<��<��<ޚ�<��<���<՚�<���<��<ۚ�<`   `   ���<��<ߚ�<S��<D��<��<��<��<K��<S��<Қ�<��<��<��<��<��<���<՚�<��<՚�<���<��<#��<��<`   `   ��<"��<1��<ޚ�<֚�<@��<)��<���<��<E��<��<��<��<&��<њ�<��<*��<Ӛ�<��<:��<��<Ś�<&��<��<`   `   ߚ�<���<���<���<��<���<4��<���<ؚ�<���<��<��<��<њ�<њ�<ʚ�<��<��<��<ʚ�<��<њ�<��<��<`   `   ˚�<���<���<1��<Ě�<���<��<��<њ�<���<��<��<��<��<ʚ�<���<��< ��<���<���<��<��<��<���<`   `   ��<��<���<���<:��<���<���<��<��<��<ޚ�<��<���<*��<��<��<���<��<���<*��<Ě�<��<ך�<��<`   `   ۚ�<+��<%��<��<��<9��<��<К�<ך�<Ț�<Ϛ�<ޚ�<՚�<Ӛ�<��< ��<��<ښ�<��<ؚ�<՚�<֚�<Ț�<ƚ�<`   `   ���<���<`��<��<3��<���<Ϛ�<��<,��<��<��<��<��<��<��<���<���<��<���<��<��<��<>��<��<`   `   ��<��<��<(��< ��<ޚ�<���<���<��<���<��<���<՚�<:��<ʚ�<���<*��<ؚ�<��<&��<��<���<���<��<`   `   [��<���<���<���<N��<$��<���<��<��<��<��<՚�<���<��<��<��<Ě�<՚�<��<��<���<��<���<$��<`   `   ���<,��<��<���< ��<��<���<��<��<ݚ�<Ϛ�<���<��<Ś�<њ�<��<��<֚�<��<���<��<��<��<��<`   `   ɚ�<0��<��<���<"��<��<���<���<<��<Ț�<Κ�<��<#��<&��<��<��<ך�<Ț�<>��<���<���<��<;��<���<`   `   ۚ�<К�<��<���< ��<-��<���<ݚ�<ך�<��<��<ۚ�<��<��<��<���<��<ƚ�<��<��<$��<��<���<-��<`   `   ���<a��<4��<)��<R��<5��<{��<+��<A��<K��<x��<]��<5��<]��<g��<K��<^��<+��<Z��<5��<o��<)��<#��<a��<`   `   a��<J��<h��<v��<��<��<���<y��<T��<��<r��<a��<_��<y��<���<D��<k��<���<+��<	��<o��<z��<I��<V��<`   `   4��<h��<#��<@��<>��<8��<$��<V��<]��<��<��<o��<ޘ�<��<c��<V��<��<8��<G��<@��<��<h��<?��<���<`   `   )��<v��<@��<&��<��<R��<d��<A��<��<���<k��<r��<���<��<J��<y��<D��<���<3��<R��<o��<��<H��<I��<`   `   R��<��<>��<��<s��<O��<���<��<h��<J��<���<J��<z��<��<f��<O��<���<��<��<��<c��<��<d��<��<`   `   5��<��<8��<R��<O��<��<P��<(��<��<6��</��<���<&��<e��<��<9��<D��<J��<+��<*��<U��<[��<Z��<\��<`   `   {��<���<$��<d��<���<P��<ܘ�<\��<3��<��<J��<\��<Ș�<P��<���<d��<��<���<y��<���<V��<s��<P��<���<`   `   +��<y��<V��<A��<��<(��<\��<���<>��<.��<���<q��<&��<i��<J��<h��<k��< ��<L��<a��<7��<>��<`��<@��<`   `   A��<T��<]��<��<h��<��<3��<>��<r��<>��<%��<��<���<��<B��<T��<X��<Y��<k��<1��<4��<1��<y��<Y��<`   `   K��<��<��<���<J��<6��<��<.��<>��<(��</��<4��<���<1��<���<A��<���<���<?��<~��<v��<2��<��<���<`   `   x��<r��<��<k��<���</��<J��<���<%��</��<���<k��<Ә�<r��<y��<I��<_��<V��<H��<B��<\��<V��<S��<I��<`   `   ]��<a��<o��<r��<J��<���<\��<q��<��<4��<k��<���<_��<S��<7��<L��<���<���<��<��<���<���<K��<-��<`   `   5��<_��<ޘ�<���<z��<&��<Ș�<&��<���<���<Ә�<_��<B��<#��<L��<]��<X��<y��<���<y��<R��<]��<V��<#��<`   `   ]��<y��<��<��<��<e��<P��<i��<��<1��<r��<S��<#��<V��<���<J��<L��<c��<o��<Z��<B��<v��<U��<%��<`   `   g��<���<c��<J��<f��<��<���<J��<B��<���<y��<7��<L��<���<{��<]��<���<?��<m��<]��<���<���<K��<7��<`   `   K��<D��<V��<y��<O��<9��<d��<h��<T��<A��<I��<L��<]��<J��<]��<���<u��<���<���<T��<B��<_��<K��<Q��<`   `   ^��<k��<��<D��<���<D��<��<k��<X��<���<_��<���<X��<L��<���<u��<��<u��<���<L��<]��<���<Y��<���<`   `   +��<���<8��<���<��<J��<���< ��<Y��<���<V��<���<y��<c��<?��<���<u��<6��<o��<{��<���<]��<��<I��<`   `   Z��<+��<G��<3��<��<+��<y��<L��<k��<?��<H��<��<���<o��<m��<���<���<o��<v��<��<H��<?��<|��<L��<`   `   5��<	��<@��<R��<��<*��<���<a��<1��<~��<B��<��<y��<Z��<]��<T��<L��<{��<��<I��<v��<"��<`��<���<`   `   o��<o��<��<o��<c��<U��<V��<7��<4��<v��<\��<���<R��<B��<���<B��<]��<���<H��<v��<K��<7��<B��<U��<`   `   )��<z��<h��<��<��<[��<s��<>��<1��<2��<V��<���<]��<v��<���<_��<���<]��<?��<"��<7��<���<Z��<��<`   `   #��<I��<?��<H��<d��<Z��<P��<`��<y��<��<S��<K��<V��<U��<K��<K��<Y��<��<|��<`��<B��<Z��<{��<H��<`   `   a��<V��<���<I��<��<\��<���<@��<Y��<���<I��<-��<#��<%��<7��<Q��<���<I��<L��<���<U��<��<H��<���<`   `   ���<���<���<��<�<���<֗�<���<���<���<���<���<���<���<���<���<Ɨ�<���<���<���<ٗ�<��<���<���<`   `   ���<���<���<ӗ�<���<ė�<���<���<���<}��<���<���<���<���<���<���<���<Ɨ�<Η�<���<Η�<ŗ�<���<���<`   `   ���<���<Y��<ʗ�<���<×�<o��<���<��<��<ؗ�<���<ӗ�<��<��<���<h��<×�< ��<ʗ�<O��<���<���<���<`   `   ��<ӗ�<ʗ�<֗�<���<՗�<���<k��<җ�<���<���<���<ߗ�<Ɨ�<r��<×�<˗�<���<ߗ�<ؗ�<Η�<��<���<���<`   `   �<���<���<���<ϗ�<���<���<���<��<z��<���<z��<���<���<t��<���<��<���<���<���<З�<���<ȗ�<���<`   `   ���<ė�<×�<՗�<���<���<ܗ�<��<���<���<���<���<��<��<���<���<˗�<ї�<Η�<���<���<���<���<���<`   `   ֗�<���<o��<���<���<ܗ�<ʗ�<ŗ�<���<��<���<ŗ�<���<ܗ�<���<���<k��<���<՗�<���<���<З�<���<���<`   `   ���<���<���<k��<���<��<ŗ�<���<���<���<���<֗�<��<{��<r��<͗�<���<���<���<���<֗�<ۗ�<���<���<`   `   ���<���<��<җ�<��<���<���<���<՗�<���<���<���<���<җ�<̗�<���<�<���<���<���<՗�<���<���<���<`   `   ���<}��<��<���<z��<���<��<���<���<��<���<h��<ߗ�<��<���<{��<���<���<���<×�<���<���<���<���<`   `   ���<���<ؗ�<���<���<���<���<���<���<���<���<���<˗�<���<���<���<_��<���<���<���<���<���<W��<���<`   `   ���<���<���<���<z��<���<ŗ�<֗�<���<h��<���<��<���<���<��<���<���<���<���<���<���<���<���<��<`   `   ���<���<ӗ�<ߗ�<���<��<���<��<���<ߗ�<˗�<���<���<��<���<���<���<���<ʗ�<���<���<���<���<��<`   `   ���<���<��<Ɨ�<���<��<ܗ�<{��<җ�<��<���<���<��<���<���<���<���<���<���<���<���<���<���<��<`   `   ���<���<��<r��<t��<���<���<r��<̗�<���<���<��<���<���<ė�<���<���<���<���<���<З�<���<���<��<`   `   ���<���<���<×�<���<���<���<͗�<���<{��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   Ɨ�<���<h��<˗�<��<˗�<k��<���<�<���<_��<���<���<���<���<���<���<���<���<���<���<���<Z��<���<`   `   ���<Ɨ�<×�<���<���<ї�<���<���<���<���<���<���<���<���<���<���<���<z��<���<���<���<���<���<���<`   `   ���<Η�< ��<ߗ�<���<Η�<՗�<���<���<���<���<���<ʗ�<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<ʗ�<ؗ�<���<���<���<���<���<×�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   ٗ�<Η�<O��<Η�<З�<���<���<֗�<՗�<���<���<���<���<���<З�<���<���<���<���<���<��<֗�<y��<���<`   `   ��<ŗ�<���<��<���<���<З�<ۗ�<���<���<���<���<���<���<���<���<���<���<���<���<֗�<���<���<���<`   `   ���<���<���<���<ȗ�<���<���<���<���<���<W��<���<���<���<���<���<Z��<���<���<���<y��<���<ۗ�<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<��<��<��<��<���<���<���<���<���<���<���<���<���<`   `   ?��<4��<;��<���<&��<3��<��<L��<U��<]��<U��<��<=��<��<L��<]��<d��<L��<
��<3��<5��<���<2��<4��<`   `   4��<b��<:��<��<��<��<��<8��< ��<���<2��<��<��<7��<��<��<2��<��<��<���<��<D��<a��<.��<`   `   ;��<:��<$��<4��<��<=��<��<Y��<��<"��<)��<���<%��<"��<��<Y��<��<=��<��<4��<��<:��<B��<+��<`   `   ���<��<4��<��<��<E��<p��<G��<��<,��<��<��<,��<���<K��<|��<>��< ��<��<>��<��<���<��<��<`   `   &��<��<��<��<��<��<N��<��<-��<��<'��<��<7��<��<>��<��<���<��<��<��</��<)��<&��<)��<`   `   3��<��<=��<E��<��<L��<��<��<0��<��<��<(��<��<'��<P��<��<>��<G��<��<-��<p��<<��<;��<t��<`   `   ��<��<��<p��<N��<��<��<.��<���<��<��<.��<ܕ�<��<U��<p��<��<��<��<D��<'��<���<$��<D��<`   `   L��<8��<Y��<G��<��<��<.��<��</��<&��<��<:��<��<��<K��<c��<2��<F��<?��<M��<$��<'��<L��<9��<`   `   U��< ��<��<��<-��<0��<���</��<���</��<��<0��<:��<��<��< ��<a��<5��<h��<'��<��<'��<o��<5��<`   `   ]��<���<"��<,��<��<��<��<&��</��<��<��<��<,��<,��<��<W��<!��<F��<B��<���<���<<��<E��<'��<`   `   U��<2��<)��<��<'��<��<��<��<��<��<7��<��<��<2��<W��<^��<>��<[��<&��<G��</��<[��<8��<^��<`   `   ��<��<���<��<��<(��<.��<:��<0��<��<��<��<��<��<���<;��<C��<��<Q��<K��<	��<J��<:��<���<`   `   =��<��<%��<,��<7��<��<ܕ�<��<:��<,��<��<��<D��<��<��<O��<'��<!��<:��<!��<$��<O��<$��<��<`   `   ��<7��<"��<���<��<'��<��<��<��<,��<2��<��<��<J��<6��<c��<���<5��<;��<���<`��<1��<I��<��<`   `   L��<��<��<K��<>��<P��<U��<K��<��<��<W��<���<��<6��<��<4��<f��<l��<Y��<4��<"��<6��<��<���<`   `   ]��<��<Y��<|��<��<��<p��<c��< ��<W��<^��<;��<O��<c��<4��<��<D��<K��<��<0��<`��<O��<:��<b��<`   `   d��<2��<��<>��<���<>��<��<2��<a��<!��<>��<C��<'��<���<f��<D��<7��<D��<d��<���<*��<C��<:��<!��<`   `   L��<��<=��< ��<��<G��<��<F��<5��<F��<[��<��<!��<5��<l��<K��<D��<h��<;��<!��<	��<_��<E��<,��<`   `   
��<��<��<��<��<��<��<?��<h��<B��<&��<Q��<:��<;��<Y��<��<d��<;��<3��<Q��<%��<B��<r��<?��<`   `   3��<���<4��<>��<��<-��<D��<M��<'��<���<G��<K��<!��<���<4��<0��<���<!��<Q��<K��<���<��<L��<O��<`   `   5��<��<��<��</��<p��<'��<$��<��<���</��<	��<$��<`��<"��<`��<*��<	��<%��<���<��<$��<��<p��<`   `   ���<D��<:��<���<)��<<��<���<'��<'��<<��<[��<J��<O��<1��<6��<O��<C��<_��<B��<��<$��<	��<;��<��<`   `   2��<a��<B��<��<&��<;��<$��<L��<o��<E��<8��<:��<$��<I��<��<:��<:��<E��<r��<L��<��<;��<3��<��<`   `   4��<.��<+��<��<)��<t��<D��<9��<5��<'��<^��<���<��<��<���<b��<!��<,��<?��<O��<p��<��<��<4��<`   `   ���<���<���<���<���<���<���<Ô�<���<���<Ҕ�<���<ߔ�<���<Δ�<���<���<Ô�<���<���<���<���<���<���<`   `   ���<���<���<���<ʔ�<Ɣ�<ܔ�<���<���<Ɣ�<��<ה�<֔�<��<Ȕ�<���<���<��<Ȕ�<Ĕ�<���<���<���<���<`   `   ���<���<ؔ�<���<���<Ҕ�<y��<���<���<���<���<���<���<���<���<���<v��<Ҕ�<���<���<Ԕ�<���<���<Ԕ�<`   `   ���<���<���<���<���<ǔ�<q��<ϔ�<���<���<��<��<���<���<є�<v��<Ĕ�<ڔ�<���<��<���<���<۔�<ܔ�<`   `   ���<ʔ�<���<���<���<���<���<֔�<ǔ�<Ô�<��<Ô�<˔�<֔�<���<���<��<���<���<ʔ�<���<���<���<���<`   `   ���<Ɣ�<Ҕ�<ǔ�<���<Ҕ�<���<ɔ�<���<���<���<���<ɔ�<���<Ԕ�<���<Ĕ�<֔�<Ȕ�<���<���<���<���<���<`   `   ���<ܔ�<y��<q��<���<���<���<ٔ�<Ô�<���<ɔ�<ٔ�<���<���<���<q��<w��<ܔ�<���<���<���<���<���<���<`   `   Ô�<���<���<ϔ�<֔�<ɔ�<ٔ�<��<���<���<��<ޔ�<ɔ�<є�<є�<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<ǔ�<���<Ô�<���<P��<���<���<���<͔�<���<���<���<���<~��<���<���<��<���<���<~��<`   `   ���<Ɣ�<���<���<Ô�<���<���<���<���<���<���<���<���<���<Ȕ�<���<v��<���<���<��<��<���<���<y��<`   `   Ҕ�<��<���<��<��<���<ɔ�<��<���<���<��<��<���<��<Ҕ�<���<���<���<���<���<���<���<���<���<`   `   ���<ה�<���<��<Ô�<���<ٔ�<ޔ�<���<���<��<���<֔�<���<o��<���<���<���<���<���<���<���<���<m��<`   `   ߔ�<֔�<���<���<˔�<ɔ�<���<ɔ�<͔�<���<���<֔�<��<���<�<���<���<Ɣ�<���<Ɣ�<���<���<Ĕ�<���<`   `   ���<��<���<���<֔�<���<���<є�<���<���<��<���<���<��<���<|��<���<i��<k��<���<{��<���<��<���<`   `   Δ�<Ȕ�<���<є�<���<Ԕ�<���<є�<���<Ȕ�<Ҕ�<o��<�<���<���<���<���<���<���<���<���<���<�<o��<`   `   ���<���<���<v��<���<���<q��<���<���<���<���<���<���<|��<���<���<���<���<���<���<{��<���<���<���<`   `   ���<���<v��<Ĕ�<��<Ĕ�<w��<���<���<v��<���<���<���<���<���<���<v��<���<���<���<���<���<���<v��<`   `   Ô�<��<Ҕ�<ڔ�<���<֔�<ܔ�<���<~��<���<���<���<Ɣ�<i��<���<���<���<���<k��<Ɣ�<���<���<���<z��<`   `   ���<Ȕ�<���<���<���<Ȕ�<���<���<���<���<���<���<���<k��<���<���<���<k��<���<���<���<���<���<���<`   `   ���<Ĕ�<���<��<ʔ�<���<���<���<���<��<���<���<Ɣ�<���<���<���<���<Ɣ�<���<���<��<���<���<���<`   `   ���<���<Ԕ�<���<���<���<���<���<��<��<���<���<���<{��<���<{��<���<���<���<��<��<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<۔�<���<���<���<���<���<���<���<���<Ĕ�<��<�<���<���<���<���<���<���<���<���<۔�<`   `   ���<���<Ԕ�<ܔ�<���<���<���<���<~��<y��<���<m��<���<���<o��<���<v��<z��<���<���<���<���<۔�<ؔ�<`   `   ���<\��<Q��<��<^��<Y��<G��<A��<a��<A��<%��<>��</��<>��<&��<A��<_��<A��<I��<Y��<\��<��<R��<\��<`   `   \��<P��<`��<5��<F��<@��<I��<f��<g��</��<��<%��<%��<��</��<h��<g��<G��<?��<H��<6��<^��<Q��<]��<`   `   Q��<`��<���<-��<<��<'��<r��<p��<k��<f��<g��<S��<h��<f��<k��<p��<r��<'��<;��<-��<���<`��<P��<��<`   `   ��<5��<-��<x��<��<F��<Y��<3��<\��<`��<.��<.��<`��<]��<3��<W��<G��<��<x��<,��<6��<��<4��<3��<`   `   ^��<F��<<��<��<-��<l��<��<,��<K��<"��<��<"��<J��<,��<��<l��<+��<��<=��<F��<]��<K��<J��<K��<`   `   Y��<@��<'��<F��<l��<B��<F��<]��<6��<S��<S��<7��<]��<E��<B��<n��<G��<&��<?��<Y��<.��<Z��<Z��<.��<`   `   G��<I��<r��<Y��<��<F��<p��<��<B��<���<@��<��<r��<F��<��<Y��<r��<I��<F��<Z��<a��<j��<a��<Z��<`   `   A��<f��<p��<3��<,��<]��<��< ��<X��<Y��< ��<��<]��<-��<3��<o��<g��<A��<n��<��<:��<:��<��<o��<`   `   a��<g��<k��<\��<K��<6��<B��<X��<6��<X��<C��<6��<J��<\��<m��<g��<`��<���<x��<0��<!��<0��<w��<���<`   `   A��</��<f��<`��<"��<S��<���<Y��<X��<���<S��<$��<`��<d��</��<B��<���<���<J��<c��<c��<J��<���<���<`   `   %��<��<g��<.��<��<S��<@��< ��<C��<S��<��<.��<h��<��<$��<^��<C��<H��<S��<5��<S��<H��<C��<^��<`   `   >��<%��<S��<.��<"��<7��<��<��<6��<$��<.��<R��<%��<?��<���<j��<(��<~��<-��<-��<~��<(��<j��<���<`   `   /��<%��<h��<`��<J��<]��<r��<]��<J��<`��<h��<%��<.��<^��<y��<e��<l��<���<t��<���<m��<e��<x��<^��<`   `   >��<��<f��<]��<,��<E��<F��<-��<\��<d��<��<?��<^��<���<C��<l��<;��<���<���<;��<l��<C��<���<^��<`   `   &��</��<k��<3��<��<B��<��<3��<m��</��<$��<���<y��<C��<���<n��<I��<���<J��<n��<���<C��<x��<���<`   `   A��<h��<p��<W��<l��<n��<Y��<o��<g��<B��<^��<j��<e��<l��<n��<^��<f��<e��<]��<o��<l��<e��<j��<]��<`   `   _��<g��<r��<G��<+��<G��<r��<g��<`��<���<C��<(��<l��<;��<I��<f��<N��<f��<I��<;��<l��<(��<C��<���<`   `   A��<G��<'��<��<��<&��<I��<A��<���<���<H��<~��<���<���<���<e��<f��<���<���<���<~��<G��<���<���<`   `   I��<?��<;��<x��<=��<?��<F��<n��<x��<J��<S��<-��<t��<���<J��<]��<I��<���<t��<-��<T��<J��<v��<n��<`   `   Y��<H��<-��<,��<F��<Y��<Z��<��<0��<c��<5��<-��<���<;��<n��<o��<;��<���<-��<5��<c��<1��<��<Y��<`   `   \��<6��<���<6��<]��<.��<a��<:��<!��<c��<S��<~��<m��<l��<���<l��<l��<~��<T��<c��< ��<:��<b��<.��<`   `   ��<^��<`��<��<K��<Z��<j��<:��<0��<J��<H��<(��<e��<C��<C��<e��<(��<G��<J��<1��<:��<h��<Z��<M��<`   `   R��<Q��<P��<4��<J��<Z��<a��<��<w��<���<C��<j��<x��<���<x��<j��<C��<���<v��<��<b��<Z��<I��<4��<`   `   \��<]��<��<3��<K��<.��<Z��<o��<���<���<^��<���<^��<^��<���<]��<���<���<n��<Y��<.��<M��<4��<��<`   `   ���<���<���<��<��<��<��<ݑ�<��<��<��<��<��<��<��<��<��<ݑ�<��<��<��<��< ��<���<`   `   ���<���<��<���<��<��<��<ϑ�<���<��<��<��<��<��<��<���<ӑ�<��<��<���<���<��<���<���<`   `   ���<��<0��<��<��<��<��<ґ�<Б�<��<��<��<��<��<͑�<ґ�<��<��<��<��<5��<��<���<��<`   `   ��<���<��<C��<��<���<%��<��<��<���<���<���<���<��< ��<��<��<��<?��<���<���<��<��<��<`   `   ��<��<��<��<ő�<��<"��<	��<��<4��<��<4��<��<	��<-��<��<���<��<$��<��<��<��<��<��<`   `   ��<��<��<���<��<��<���<��<(��<��<��<.��<��<���<��<��<��<��<��<��<��<���<���< ��<`   `   ��<��<��<%��<"��<���<��<!��< ��<���<���<!��<$��<���<��<%��<��<��<��<���<��<ґ�<��<���<`   `   ݑ�<ϑ�<ґ�<��<	��<��<!��<"��<���< ��<&��<��<��<��< ��<ˑ�<ӑ�<��<ܑ�<��<��<��<��<���<`   `   ��<���<Б�<��<��<(��< ��<���<:��<���<��<(��<��<��<ّ�<���<��<Ñ�<Ǒ�<��<��<��<�<Ñ�<`   `   ��<��<��<���<4��<��<���< ��<���<���<��<<��<���<ߑ�<��<��<��<ɑ�<��<ޑ�<���<��<ʑ�<��<`   `   ��<��<��<���<��<��<���<&��<��<��<��<���<��<��<��<��<��<���<!��<��<��<���<���<��<`   `   ��<��<��<���<4��<.��<!��<��<(��<<��<���<��<��<!��<��<Ց�<���<��<��<
��<��<��<֑�<��<`   `   ��<��<��<���<��<��<$��<��<��<���<��<��<��<���<Б�<���<��<���<���<���<��<���<͑�<���<`   `   ��<��<��<��<	��<���<���<��<��<ߑ�<��<!��<���<��<��<���<��<��<��<��<���<��<��<���<`   `   ��<��<͑�< ��<-��<��<��< ��<ّ�<��<��<��<Б�<��<֑�<ё�<��<��<���<ё�<ё�<��<Б�<��<`   `   ��<���<ґ�<��<��<��<%��<ˑ�<���<��<��<Ց�<���<���<ё�<��<��<ݑ�<��<ӑ�<���<���<֑�<ߑ�<`   `   ��<ӑ�<��<��<���<��<��<ӑ�<��<��<��<���<��<��<��<��<��<��<��<��<��<���<���<��<`   `   ݑ�<��<��<��<��<��<��<��<Ñ�<ɑ�<���<��<���<��<��<ݑ�<��<��<��<���<��<��<ʑ�<ɑ�<`   `   ��<��<��<?��<$��<��<��<ܑ�<Ǒ�<��<!��<��<���<��<���<��<��<��<���<��<"��<��<���<ܑ�<`   `   ��<���<��<���<��<��<���<��<��<ޑ�<��<
��<���<��<ё�<ӑ�<��<���<��<��<���<��<��<���<`   `   ��<���<5��<���<��<��<��<��<��<���<��<��<��<���<ё�<���<��<��<"��<���<���<��<��<��<`   `   ��<��<��<��<��<���<ґ�<��<��<��<���<��<���<��<��<���<���<��<��<��<��<ʑ�<���<��<`   `    ��<���<���<��<��<���<��<��<�<ʑ�<���<֑�<͑�<��<Б�<֑�<���<ʑ�<���<��<��<���<��<��<`   `   ���<���<��<��<��< ��<���<���<Ñ�<��<��<��<���<���<��<ߑ�<��<ɑ�<ܑ�<���<��<��<��<��<`   `   r��<֐�<���<���<���<���<���<
��<А�<���<���<���<���<���<���<���<���<
��<Ԑ�<���<���<���<���<֐�<`   `   ֐�<���<���<ؐ�<̐�<���<���<ϐ�<Ӑ�<ߐ�<���<���<���<���<ڐ�<ސ�<א�<���<���<ڐ�<ܐ�<}��<���<ݐ�<`   `   ���<���<���<���<���<���<�<���<А�<���<���<���<���<���<ː�<���<Ȑ�<���<���<���<���<���<���<��<`   `   ���<ؐ�<���<W��<Ր�<���<o��<֐�<��<���<���<���<���<��<ѐ�<b��<���<��<P��<~��<ܐ�<���<͐�<ː�<`   `   ���<̐�<���<Ր�<���<���<���<���<���<���<���<���<���<���<���<���<ߐ�<Ր�<���<̐�<���<А�<���<А�<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<͐�<���<���<ɐ�<`   `   ���<���<�<o��<���<���<���<���<Ґ�<���<Ð�<���<���<���<���<o��<Ɛ�<���<���<���<ϐ�<���<Ґ�<���<`   `   
��<ϐ�<���<֐�<���<���<���<ϐ�<���<Ð�<Ԑ�<���<���<��<ѐ�<���<א�<��<ߐ�<���<ɐ�<Ɛ�<���<��<`   `   А�<Ӑ�<А�<��<���<���<Ґ�<���<���<���<ې�<���<���<��<��<Ӑ�<���<��<Ȑ�<��<Ґ�<��<���<��<`   `   ���<ߐ�<���<���<���<���<���<Ð�<���<���<���<ϐ�<���<���<ڐ�<���<���<���<ސ�<���<���<��<���<���<`   `   ���<���<���<���<���<���<Ð�<Ԑ�<ې�<���<���<���<���<���<���<���<
��<���<���<���<���<���<��<���<`   `   ���<���<���<���<���<���<���<���<���<ϐ�<���<���<���<���<���<Ր�<��<���<���<��<���<��<א�<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<А�<Ð�<��<Ð�<Ԑ�<���<���<���<`   `   ���<���<���<��<���<���<���<��<��<���<���<���<���<-��<��<���<��<��<��<���<���<��<.��<���<`   `   ���<ڐ�<ː�<ѐ�<���<���<���<ѐ�<��<ڐ�<���<���<���<��<���<ߐ�<��<���<��<ߐ�<���<��<���<���<`   `   ���<ސ�<���<b��<���<���<o��<���<Ӑ�<���<���<Ր�<���<���<ߐ�<���<���<���<���<��<���<���<א�<���<`   `   ���<א�<Ȑ�<���<ߐ�<���<Ɛ�<א�<���<���<
��<��<А�<��<��<���<��<���<��<��<͐�<��<��<���<`   `   
��<���<���<��<Ր�<���<���<��<��<���<���<���<Ð�<��<���<���<���<���<��<�<���<���<���<���<`   `   Ԑ�<���<���<P��<���<���<���<ߐ�<Ȑ�<ސ�<���<���<��<��<��<���<��<��<��<���<���<ސ�<���<ߐ�<`   `   ���<ڐ�<���<~��<̐�<���<���<���<��<���<���<��<Ð�<���<ߐ�<��<��<�<���<���<���<���<���<���<`   `   ���<ܐ�<���<ܐ�<���<͐�<ϐ�<ɐ�<Ґ�<���<���<���<Ԑ�<���<���<���<͐�<���<���<���<Đ�<ɐ�<ې�<͐�<`   `   ���<}��<���<���<А�<���<���<Ɛ�<��<��<���<��<���<��<��<���<��<���<ސ�<���<ɐ�<���<���<ސ�<`   `   ���<���<���<͐�<���<���<Ґ�<���<���<���<��<א�<���<.��<���<א�<��<���<���<���<ې�<���<���<͐�<`   `   ֐�<ݐ�<��<ː�<А�<ɐ�<���<��<��<���<���<���<���<���<���<���<���<���<ߐ�<���<͐�<ސ�<͐�<ې�<`   `   ���<���<���<���<m��<���<`��<>��<c��<~��<y��<���<���<���<���<~��<J��<>��<|��<���<U��<���<���<���<`   `   ���<֏�<���<~��<���<���<W��<p��<���<���<���<���<���<|��<}��<���<{��<D��<���<̏�<���<x��<؏�<���<`   `   ���<���<���<���<���<p��<���<���<l��<���<���<���<���<���<f��<���<���<p��<���<���<���<���<���<��<`   `   ���<~��<���<Ǐ�<���<b��<���<o��<~��<���<���<���<���<���<h��<���<m��<���<���<���<���<ď�<���<���<`   `   m��<���<���<���<���<я�<r��<~��<{��<���<r��<���<l��<~��<���<я�<e��<���<ʏ�<���<^��<���<b��<���<`   `   ���<���<p��<b��<я�<���<���<���<���<���<���<���<���<{��<���<��<m��<`��<���<���<���<u��<w��<���<`   `   `��<W��<���<���<r��<���<���<���<���<��<���<���<��<���<g��<���<���<W��<a��<���<Џ�<���<ԏ�<���<`   `   >��<p��<���<o��<~��<���<���<+��<���<���<2��<n��<���<���<h��<���<{��<H��<���<p��<W��<Q��<r��<���<`   `   c��<���<l��<~��<{��<���<���<���<Q��<���<���<���<g��<~��<���<���<N��<���<u��<{��<f��<{��<j��<���<`   `   ~��<���<���<���<���<���<��<���<���<Џ�<���<���<���<z��<}��<���<���<p��<���<���<���<���<q��<��<`   `   y��<���<���<���<r��<���<���<2��<���<���<X��<���<Ï�<���<w��<���<i��<c��<���<���<���<c��<r��<���<`   `   ���<���<���<���<���<���<���<n��<���<���<���<���<���<���<͏�<���<p��<���<r��<|��<���<e��<���<Տ�<`   `   ���<���<���<���<l��<���<��<���<g��<���<Ï�<���<~��<x��<r��<d��<���<l��<H��<l��<���<d��<i��<x��<`   `   ���<|��<���<���<~��<{��<���<���<~��<z��<���<���<x��<J��<s��<���<R��<���<}��<G��<���<{��<L��<w��<`   `   ���<}��<f��<h��<���<���<g��<h��<���<}��<w��<͏�<r��<s��<���<y��<M��<���<b��<y��<���<s��<r��<͏�<`   `   ~��<���<���<���<я�<��<���<���<���<���<���<���<d��<���<y��<i��<~��<s��<_��<���<���<b��<���<���<`   `   J��<{��<���<m��<e��<m��<���<{��<N��<���<i��<p��<���<R��<M��<~��<���<~��<O��<R��<���<p��<n��<���<`   `   >��<D��<p��<���<���<`��<W��<H��<���<p��<c��<���<l��<���<���<s��<~��<���<}��<j��<���<\��<q��<���<`   `   |��<���<���<���<ʏ�<���<a��<���<u��<���<���<r��<H��<}��<b��<_��<O��<}��<S��<r��<���<���<f��<���<`   `   ���<̏�<���<���<���<���<���<p��<{��<���<���<|��<l��<G��<y��<���<R��<j��<r��<z��<���<���<r��<���<`   `   U��<���<���<���<^��<���<Џ�<W��<f��<���<���<���<���<���<���<���<���<���<���<���<S��<W��<���<���<`   `   ���<x��<���<ď�<���<u��<���<Q��<{��<���<c��<e��<d��<{��<s��<b��<p��<\��<���<���<W��<���<w��<���<`   `   ���<؏�<���<���<b��<w��<ԏ�<r��<j��<q��<r��<���<i��<L��<r��<���<n��<q��<f��<r��<���<w��<N��<���<`   `   ���<���<��<���<���<���<���<���<���<��<���<Տ�<x��<w��<͏�<���<���<���<���<���<���<���<���<��<`   `   P��<s��<{��<|��<P��<���<���<���<���<���<8��<b��<l��<b��<J��<���<���<���<���<���<3��<|��<���<s��<`   `   s��<S��<V��<N��<b��<���<���<M��<���<���<e��<e��<g��<^��<���<���<[��<v��<���<x��<U��<D��<T��<}��<`   `   {��<V��<���<O��<2��<Q��<���<:��<W��<~��<j��<��<o��<~��<R��<:��<���<Q��<)��<O��<���<V��<p��<r��<`   `   |��<N��<O��<���<���<2��<`��<���<���<[��<W��<P��<]��<���<���<K��<@��<���<���<=��<U��<���<���<���<`   `   P��<b��<2��<���<D��<m��<t��<���<I��<���<���<���<6��<���<���<m��< ��<���<R��<b��<>��<���<~��<���<`   `   ���<���<Q��<2��<m��<p��<*��<`��<���<>��<E��<���<c��<��<f��<���<@��<?��<���<���<M��<k��<l��<F��<`   `   ���<���<���<`��<t��<*��<h��<g��<q��<��<Z��<g��<{��<*��<h��<`��<���<���<���<]��<s��<Z��<z��<]��<`   `   ���<M��<:��<���<���<`��<g��<v��<���<���<}��<R��<c��<���<���<'��<[��<���<���<���<���<���<���<���<`   `   ���<���<W��<���<I��<���<q��<���<M��<���<��<���<0��<���<t��<���<���<���<J��<���<���<���<<��<���<`   `   ���<���<~��<[��<���<>��<��<���<���<���<E��<���<]��<l��<���<Ď�<���<~��<h��<_��<g��<u��<��<���<`   `   8��<e��<j��<W��<���<E��<Z��<}��<��<E��<~��<W��<z��<e��<8��<I��<���<���<���<`��<l��<���<���<I��<`   `   b��<e��<��<P��<���<���<g��<R��<���<���<W��<	��<g��<m��<��<f��<n��<���<���<���<���<`��<g��<���<`   `   l��<g��<o��<]��<6��<c��<{��<c��<0��<]��<z��<g��<_��<|��<���<���<���<���<p��<���<���<���<���<|��<`   `   b��<^��<~��<���<���<��<*��<���<���<l��<e��<m��<|��<t��<���<z��<S��<���<���<E��<���<���<u��<z��<`   `   J��<���<R��<���<���<f��<h��<���<t��<���<8��<��<���<���<���<���<t��<ǎ�<���<���<��<���<���<��<`   `   ���<���<:��<K��<m��<���<`��<(��<���<Ď�<I��<f��<���<z��<���<���<y��<k��<���<���<���<���<g��<A��<`   `   ���<[��<���<@��< ��<@��<���<[��<���<���<���<n��<���<S��<t��<y��<J��<y��<w��<S��<���<n��<���<���<`   `   ���<v��<Q��<���<���<?��<���<���<���<~��<���<���<���<���<ǎ�<k��<y��<Ҏ�<���<���<���<���<��<���<`   `   ���<���<)��<���<R��<���<���<���<J��<h��<���<���<p��<���<���<���<w��<���<���<���<���<h��<:��<���<`   `   ���<x��<O��<=��<b��<���<]��<���<���<_��<`��<���<���<E��<���<���<S��<���<���<Y��<g��<���<���<G��<`   `   3��<U��<���<U��<>��<M��<s��<���<���<g��<l��<���<���<���<��<���<���<���<���<g��<���<���<���<M��<`   `   |��<D��<V��<���<���<k��<Z��<���<���<u��<���<`��<���<���<���<���<n��<���<h��<���<���<E��<l��<���<`   `   ���<T��<p��<���<~��<l��<z��<���<<��<��<���<g��<���<u��<���<g��<���<��<:��<���<���<l��<g��<���<`   `   s��<}��<r��<���<���<F��<]��<���<���<���<I��<���<|��<z��<��<A��<���<���<���<G��<M��<���<���<`��<`   `   :��<��<y��<L��<���<���<!��<���<U��<Z��<V��<y��<m��<y��<i��<Z��<4��<���<G��<���<o��<L��<���<��<`   `   ��<C��<]��<x��<���<b��<F��<L��<m��<o��<o��<���<���<h��<c��<}��<\��</��<R��<���<���<J��<C��<���<`   `   y��<]��<ߍ�<]��< ��<b��<���<F��<S��<D��<���<|��<���<D��<O��<F��<���<b��<��<]��<��<]��<n��<���<`   `   L��<x��<]��<a��<���<w��<B��<���<���<V��<r��<k��<Y��<���<���<+��<���<���<Q��<J��<���<V��<*��<*��<`   `   ���<���< ��<���<���<w��<Q��<���<6��<|��<���<|��<"��<���<t��<w��<f��<���<C��<���<|��<k��<(��<k��<`   `   ���<b��<b��<w��<w��<���<���<b��<v��<}��<���<���<f��<o��<���<���<���<O��<R��<���<���<���<���<|��<`   `   !��<F��<���<B��<Q��<���<���<I��<���<V��<~��<I��<���<���<F��<B��<���<F��<&��<��<m��<5��<v��<��<`   `   ���<L��<F��<���<���<b��<I��<���<���<���<���<2��<f��<���<���<3��<\��<���<m��<���<M��<C��<���<|��<`   `   U��<m��<S��<���<6��<v��<���<���<��<���<���<v��<��<���<r��<m��<:��<N��<Z��<}��<Q��<}��<K��<N��<`   `   Z��<o��<D��<V��<|��<}��<V��<���<���<?��<���<���<Y��<1��<c��<d��<��<t��<`��<5��<?��<p��<t��<	��<`   `   V��<o��<���<r��<���<���<~��<���<���<���<h��<r��<���<o��<W��<W��<���<s��<V��<���<<��<s��<ō�<W��<`   `   y��<���<|��<k��<|��<���<I��<2��<v��<���<r��<i��<���<���<f��<m��<8��<��<w��<���<
��<(��<m��<r��<`   `   m��<���<���<Y��<"��<f��<���<f��<��<Y��<���<���<^��<T��<_��<O��<i��<a��<;��<a��<p��<O��<S��<T��<`   `   y��<h��<D��<���<���<o��<���<���<���<1��<o��<���<T��<_��<V��<C��<u��<[��<L��<e��<L��<b��<_��<P��<`   `   i��<c��<O��<���<t��<���<F��<���<r��<c��<W��<f��<_��<V��<��<f��</��<��<O��<f��<��<V��<c��<f��<`   `   Z��<}��<F��<+��<w��<���<B��<3��<m��<d��<W��<m��<O��<C��<f��<���<M��<<��<���<s��<L��<K��<m��<P��<`   `   4��<\��<���<���<f��<���<���<\��<:��<��<���<8��<i��<u��</��<M��<���<M��<2��<u��<c��<8��<���<��<`   `   ���</��<b��<���<���<O��<F��<���<N��<t��<s��<��<a��<[��<��<<��<M��<��<L��<^��<
��<l��<t��<^��<`   `   G��<R��<��<Q��<C��<R��<&��<m��<Z��<`��<V��<w��<;��<L��<O��<���<2��<L��<N��<w��<S��<`��<J��<m��<`   `   ���<���<]��<J��<���<���<��<���<}��<5��<���<���<a��<e��<f��<s��<u��<^��<w��<���<?��<���<���< ��<`   `   o��<���<��<���<|��<���<m��<M��<Q��<?��<<��<
��<p��<L��<��<L��<c��<
��<S��<?��<7��<M��<���<���<`   `   L��<J��<]��<V��<k��<���<5��<C��<}��<p��<s��<(��<O��<b��<V��<K��<8��<l��<`��<���<M��<��<���<���<`   `   ���<C��<n��<*��<(��<���<v��<���<K��<t��<ō�<m��<S��<_��<c��<m��<���<t��<J��<���<���<���<��<*��<`   `   ��<���<���<*��<k��<|��<��<|��<N��<	��<W��<r��<T��<P��<f��<P��<��<^��<m��< ��<���<���<*��<���<`   `   Z��<W��<���<���<5��<��<[��<���<���<���<���<���<~��<���<���<���<j��<���<���<��<��<���<���<W��<`   `   W��<���<i��<��<���<���<A��<O��<���<r��<Y��<+��<0��<S��<d��<���<b��<+��<���<���<"��<W��<���<a��<`   `   ���<i��<V��<i��<���<w��<���<���<i��<@��<���<K��<���<@��<h��<���<���<w��<���<i��<]��<i��<���<1��<`   `   ���<��<i��<���<D��<F��<d��<���<u��<���<W��<Q��<���<���<s��<N��<X��<[��<���<W��<"��<���<���<���<`   `   5��<���<���<D��<��<���<��<F��<r��<y��<��<y��<]��<F��<:��<���<��<D��<���<���<!��<���<n��<���<`   `   ��<���<w��<F��<���<���<E��<~��<���<a��<g��<���<���</��<���<���<X��<d��<���<���<^��<g��<f��<S��<`   `   [��<A��<���<d��<��<E��<Ì�<@��<l��<j��<V��<@��<Ԍ�<E��<��<d��<���<A��<c��<s��<���<T��<���<s��<`   `   ���<O��<���<���<F��<~��<@��<5��<x��<���<:��<)��<���<]��<s��<��<b��<���<���<���<n��<c��<���<���<`   `   ���<���<i��<u��<r��<���<l��<x��<)��<x��<|��<���<V��<u��<���<���<p��<���<I��<{��<���<{��<8��<���<`   `   ���<r��<@��<���<y��<a��<j��<���<x��<T��<g��<���<���<-��<d��<���<O��<k��<���<���<���<���<j��<<��<`   `   ���<Y��<���<W��<��<g��<V��<:��<|��<g��<���<W��<���<Y��<���<���<���<l��<���<���<��<l��<���<���<`   `   ���<+��<K��<Q��<y��<���<@��<)��<���<���<W��<8��<0��<���<x��<o��<j��<}��<z��<���<���<W��<n��<���<`   `   ~��<0��<���<���<]��<���<Ԍ�<���<V��<���<���<0��<o��<v��<L��<���<Č�<���<#��<���<̌�<���<@��<v��<`   `   ���<S��<@��<���<F��</��<E��<]��<u��<-��<Y��<���<v��<���<���<s��<v��<���<���<d��<~��<���<���<q��<`   `   ���<d��<h��<s��<:��<���<��<s��<���<d��<���<x��<L��<���<���<���<d��<�<���<���<���<���<S��<x��<`   `   ���<���<���<N��<���<���<d��<��<���<���<���<o��<���<s��<���<u��<t��<b��<c��<���<~��<���<n��<���<`   `   j��<b��<���<X��<��<X��<���<b��<p��<O��<���<j��<Č�<v��<d��<t��<��<t��<h��<v��<���<j��<���<O��<`   `   ���<+��<w��<[��<D��<d��<A��<���<���<k��<l��<}��<���<���<�<b��<t��<Ќ�<���<���<���<f��<j��<���<`   `   ���<���<���<���<���<���<c��<���<I��<���<���<z��<#��<���<���<c��<h��<���<:��<z��<���<���<:��<���<`   `   ��<���<i��<W��<���<���<s��<���<{��<���<���<���<���<d��<���<���<v��<���<z��<���<���<���<���<]��<`   `   ��<"��<]��<"��<!��<^��<���<n��<���<���<��<���<̌�<~��<���<~��<���<���<���<���<j��<n��<Ì�<^��<`   `   ���<W��<i��<���<���<g��<T��<c��<{��<���<l��<W��<���<���<���<���<j��<f��<���<���<n��<>��<f��<���<`   `   ���<���<���<���<n��<f��<���<���<8��<j��<���<n��<@��<���<S��<n��<���<j��<:��<���<Ì�<f��<Y��<���<`   `   W��<a��<1��<���<���<S��<s��<���<���<<��<���<���<v��<q��<x��<���<O��<���<���<]��<^��<���<���<��<`   `   ��<���<p��<���<���<���<���<���<���<���<I��<���<ċ�<���<]��<���<s��<���<���<���<j��<���<���<���<`   `   ���<���<���<���<���<���<��<@��<���<���<���<���<���<���<���<���<T��<k��<���<���<���<q��<���<���<`   `   p��<���<��<���<7��<~��<ċ�<[��<y��<���<ŋ�<���<Ë�<���<z��<[��<ċ�<~��<5��<���<��<���<j��<6��<`   `   ���<���<���<���<���<}��<t��<ċ�<���<l��<���<���<s��<���<���<`��<���<Ӌ�<���<w��<���<Ë�<���<���<`   `   ���<���<7��<���<���<���<���<Ћ�<v��<���<�<���<a��<Ћ�<���<���<~��<���<[��<���<w��<���<���<���<`   `   ���<���<~��<}��<���<Ƌ�<l��<���<���<���<���<���<���<X��<���<͋�<���<n��<���<���<j��<n��<l��<^��<`   `   ���<��<ċ�<t��<���<l��<���<���<���<g��<���<���<���<l��<���<t��<���<��<���<���<���<z��<���<���<`   `   ���<@��<[��<ċ�<Ћ�<���<���<���<���<���<ŋ�<���<���<��<���<J��<T��<���<p��<d��<���<���<a��<���<`   `   ���<���<y��<���<v��<���<���<���<p��<���<���<���<Z��<���<���<���<y��<���<P��<���<���<���<@��<���<`   `   ���<���<���<l��<���<���<g��<���<���<S��<���<���<s��<x��<���<���<���<���<���<Y��<e��<���<���<���<`   `   I��<���<ŋ�<���<Ë�<���<���<ŋ�<���<���<���<���<ϋ�<���<P��<{��<x��<c��<z��<��<[��<c��<���<{��<`   `   ���<���<���<���<���<���<���<���<���<���<���<t��<���<���<q��<���<p��<���<���<���<���<\��<���<���<`   `   ċ�<���<Ë�<s��<a��<���<���<���<Z��<s��<ϋ�<���<���<���<~��<���<���<���<V��<���<���<���<q��<���<`   `   ���<���<���<���<Ћ�<X��<l��<��<���<x��<���<���<���<���<v��<*��< ��<���<���<��<6��<���<���<���<`   `   ]��<���<z��<���<���<���<���<���<���<���<P��<q��<~��<v��<w��<���<f��<���<���<���<[��<v��<���<q��<`   `   ���<���<[��<`��<���<͋�<t��<J��<���<���<{��<���<���<*��<���<���<N��<:��<���<�<6��<���<���<w��<`   `   s��<T��<ċ�<���<~��<���<���<T��<y��<���<x��<p��<���< ��<f��<N��<���<N��<j��< ��<���<p��<��<���<`   `   ���<k��<~��<Ӌ�<���<n��<��<���<���<���<c��<���<���<���<���<:��<N��<Ë�<���<z��<���<_��<���<���<`   `   ���<���<5��<���<[��<���<���<p��<P��<���<z��<���<V��<���<���<���<j��<���<o��<���<q��<���<E��<p��<`   `   ���<���<���<w��<���<���<���<d��<���<Y��<��<���<���<��<���<�< ��<z��<���<��<e��<���<a��<v��<`   `   j��<���<��<���<w��<j��<���<���<���<e��<[��<���<���<6��<[��<6��<���<���<q��<e��<���<���<ɋ�<j��<`   `   ���<q��<���<Ë�<���<n��<z��<���<���<���<c��<\��<���<���<v��<���<p��<_��<���<���<���<f��<l��<���<`   `   ���<���<j��<���<���<l��<���<a��<@��<���<���<���<q��<���<���<���<��<���<E��<a��<ɋ�<l��<u��<���<`   `   ���<���<6��<���<���<^��<���<���<���<���<{��<���<���<���<q��<w��<���<���<p��<v��<j��<���<���<%��<`   `   ى�<���<Ȋ�<���<܊�<���<���<���<Ê�<���<���<���<���<���<���<���<���<���<���<���<���<���<ڊ�<���<`   `   ���<ϊ�<���<���<��<ڊ�<ϊ�<ъ�<��<���<Ċ�<���<���<�<���<���<��<���<Ǌ�<���<���<v��<ˊ�<Ɗ�<`   `   Ȋ�<���<��<���<q��<���<'��<���<���<���<Ŋ�<���<���<���<���<���<$��<���<r��<���<���<���<Ɗ�<��<`   `   ���<���<���<׊�<��<���<���<���<���<���<���<���<���<���<���<���<���<���<Ŋ�<���<���<���<���<���<`   `   ܊�<��<q��<��<���<���<���<ي�<���<̊�<���<̊�<���<ي�<���<���<���<��<���<��<Ɋ�<Ǌ�<���<Ǌ�<`   `   ���<ڊ�<���<���<���<���<���<���<���<���<���<Ċ�<���<���<���<���<���<���<Ǌ�<Ǌ�<���<��<��<���<`   `   ���<ϊ�<'��<���<���<���<��<���<���<���<���<���<��<���<���<���<!��<ϊ�<���<���<؊�<���<��<���<`   `   ���<ъ�<���<���<ي�<���<���<���<���<���<���<���<���<��<���<���<��<���<Ҋ�<��<���<���<��<��<`   `   Ê�<��<���<���<���<���<���<���<T��<���<ʊ�<���<���<���<���<��<���<���<���<Ҋ�<ϊ�<Ҋ�<���<���<`   `   ���<���<���<���<̊�<���<���<���<���<���<���<ފ�<���<���<���<���<���<Ɋ�<��<Ȋ�<Պ�<���<Ŋ�<���<`   `   ���<Ċ�<Ŋ�<���<���<���<���<���<ʊ�<���<���<���<̊�<Ċ�<���<ϊ�<ъ�<���<ߊ�<��<���<���<��<ϊ�<`   `   ���<���<���<���<̊�<Ċ�<���<���<���<ފ�<���<���<���<���<��<��<���<���<���<	��<���<���<���<���<`   `   ���<���<���<���<���<���<��<���<���<���<̊�<���<���<���<���<ˊ�<���<���<���<���<��<ˊ�<���<���<`   `   ���<�<���<���<ي�<���<���<��<���<���<Ċ�<���<���<�<ي�<׊�<��<���<͊�<ڊ�<��<��<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<���<��<���<ي�<���<��<���<���<͊�<��<���<ي�<Ɗ�<��<`   `   ���<���<���<���<���<���<���<���<��<���<ϊ�<��<ˊ�<׊�<��<Պ�<Ċ�<���<�<���<��<Ċ�<���<͊�<`   `   ���<��<$��<���<���<���<!��<��<���<���<ъ�<���<���<��<���<Ċ�<���<Ċ�<���<��<���<���<׊�<���<`   `   ���<���<���<���<��<���<ϊ�<���<���<Ɋ�<���<���<���<���<���<���<Ċ�<���<͊�<���<���<���<Ŋ�<���<`   `   ���<Ǌ�<r��<Ŋ�<���<Ǌ�<���<Ҋ�<���<��<ߊ�<���<���<͊�<͊�<�<���<͊�<���<���<Ԋ�<��<���<Ҋ�<`   `   ���<���<���<���<��<Ǌ�<���<��<Ҋ�<Ȋ�<��<	��<���<ڊ�<��<���<��<���<���<��<Պ�<݊�<��<���<`   `   ���<���<���<���<Ɋ�<���<؊�<���<ϊ�<Պ�<���<���<��<��<���<��<���<���<Ԋ�<Պ�<���<���<��<���<`   `   ���<v��<���<���<Ǌ�<��<���<���<Ҋ�<���<���<���<ˊ�<��<ي�<Ċ�<���<���<��<݊�<���<���<��<ي�<`   `   ڊ�<ˊ�<Ɗ�<���<���<��<��<��<���<Ŋ�<��<���<���<���<Ɗ�<���<׊�<Ŋ�<���<��<��<��<���<���<`   `   ���<Ɗ�<��<���<Ǌ�<���<���<��<���<���<ϊ�<���<���<���<��<͊�<���<���<Ҋ�<���<���<ي�<���<��<`   `   ���<���<���<��<��<ۉ�<݉�<���<*��<���<Չ�<��<���<��<��<���<��<���<���<ۉ�<׉�<��<��<���<`   `   ���<��< ��<���<��<I��<ĉ�<���<���<���<ى�<��<��<ى�<��<��<ʉ�<���<7��<��<ǉ�<��<��<��<`   `   ���< ��<!��<��<��<̉�<��<��<��<���<
��<	��<��<���<��<��<��<̉�<��<��<��< ��<���<���<`   `   ��<���<��<9��<܉�<щ�<(��<��<(��<!��<��<��<)��<0��<��<��<��<��<(��<ى�<ǉ�<
��<��<��<`   `   ��<��<��<܉�<
��<Q��<��<މ�<��<$��<���<$��<��<މ�<��<Q��<��<܉�<*��<��<��<,��<щ�<,��<`   `   ۉ�<I��<̉�<щ�<Q��</��<��<���<%��<ى�<ى�<-��<��<��<!��<_��<��<�<7��<߉�<ډ�<��<��<͉�<`   `   ݉�<ĉ�<��<(��<��<��<F��<��<��<"��<��<��<K��<��<��<(��<��<ĉ�<��<؉�<��<��<��<؉�<`   `   ���<���<��<��<މ�<���<��<ŉ�<&��<.��<ŉ�<���<��<��<��<݉�<ʉ�<���<?��<��<���<���<��<Q��<`   `   *��<���<��<(��<��<%��<��<&��<��<&��< ��<%��<���<(��<���<���<��<��<���<��<��<��<���<��<`   `   ���<���<���<!��<$��<ى�<"��<.��<&��<��<ى�<2��<)��<��<��<��<��<��<ω�<�<Ή�<���<݉�<ډ�<`   `   Չ�<ى�<
��<��<���<ى�<��<ŉ�< ��<ى�<���<��<��<ى�<��<��<��<(��<��<��<Љ�<(��</��<��<`   `   ��<��<	��<��<$��<-��<��<���<%��<2��<��<���<��<��<��<���<���<ω�<މ�<��<ۉ�<��<���<%��<`   `   ���<��<��<)��<��<��<K��<��<���<)��<��<��<���<���<���<���<!��<���<���<���<'��<���<���<���<`   `   ��<ى�<���<0��<މ�<��<��<��<(��<��<ى�<��<���<��<��<݉�<��<,��<��<���<��<'��<��<���<`   `   ��<��<��<��<��<!��<��<��<���<��<��<��<���<��<�<���<��<���<��<���<���<��<ĉ�<��<`   `   ���<��<��<��<Q��<_��<(��<݉�<���<��<��<���<���<݉�<���<��<Ή�<���<��<É�<��<���<���<��<`   `   ��<ʉ�<��<��<��<��<��<ʉ�<��<��<��<���<!��<��<��<Ή�<���<Ή�<��<��<��<���<��<��<`   `   ���<���<̉�<��<܉�<�<ĉ�<���<��<��<(��<ω�<���<,��<���<���<Ή�<��<��<���<ۉ�<(��<݉�<��<`   `   ���<7��<��<(��<*��<7��<��<?��<���<ω�<��<މ�<���<��<��<��<��<��<؉�<މ�<��<ω�<���<?��<`   `   ۉ�<��<��<ى�<��<߉�<؉�<��<��<�<��<��<���<���<���<É�<��<���<މ�<��<Ή�<��<��<ˉ�<`   `   ׉�<ǉ�<��<ǉ�<��<ډ�<��<���<��<Ή�<Љ�<ۉ�<'��<��<���<��<��<ۉ�<��<Ή�<��<���<��<ډ�<`   `   ��<��< ��<
��<,��<��<��<���<��<���<(��<��<���<'��<��<���<���<(��<ω�<��<���<׉�<��<:��<`   `   ��<��<���<��<щ�<��<��<��<���<݉�</��<���<���<��<ĉ�<���<��<݉�<���<��<��<��<ȉ�<��<`   `   ���<��<���<��<,��<͉�<؉�<Q��<��<ډ�<��<%��<���<���<��<��<��<��<?��<ˉ�<ډ�<:��<��<��<`   `   	��<O��<��<m��<[��<U��<C��<C��<r��<W��<)��<R��<M��<R��<5��<W��<]��<C��<Z��<U��<G��<m��<��<O��<`   `   O��<��<Q��<3��<1��<l��<Y��<)��<G��<v��<f��<T��<\��<h��<i��<K��<9��<P��<]��<9��<?��<K��<	��<P��<`   `   ��<Q��<���<F��<)��<Z��<���<?��<;��<D��<I��<J��<@��<D��<C��<?��<���<Z��</��<F��<���<Q��<��<���<`   `   m��<3��<F��<b��<V��<5��<*��<o��<L��<���<M��<N��<��<P��<b��<"��<E��<_��<S��<@��<?��<n��<a��<g��<`   `   [��<1��<)��<V��<p��<!��<��<b��<��<I��<k��<I��<��<b��<&��<!��<W��<V��<>��<1��<O��<l��<
��<l��<`   `   U��<l��<Z��<5��<!��<*��<V��<,��<H��<S��<R��<M��<4��<N��<��<*��<E��<T��<]��<V��<s��<H��<B��<h��<`   `   C��<Y��<���<*��<��<V��<q��<I��<T��<#��<P��<I��<r��<V��<��<*��<���<Y��<Q��<R��<e��<m��<v��<R��<`   `   C��<)��<?��<o��<b��<,��<I��<Q��<*��<.��<O��<A��<4��<k��<b��<9��<9��<D��<E��<#��<F��<;��<��<T��<`   `   r��<G��<;��<L��<��<H��<T��<*��<��<*��<]��<H��<	��<L��<N��<G��<a��<S��<6��<o��<���<o��<,��<S��<`   `   W��<v��<D��<���<I��<S��<#��<.��<*��<��<R��<R��<��<>��<i��<W��<F��<U��<���<U��<`��<���<P��<7��<`   `   )��<f��<I��<M��<k��<R��<P��<O��<]��<R��<c��<M��<H��<f��<5��<?��<=��<J��<a��<T��<F��<J��<R��<?��<`   `   R��<T��<J��<N��<I��<M��<I��<A��<H��<R��<M��<D��<\��<R��<o��<v��<Z��<E��<���<���<P��<K��<p��<|��<`   `   M��<\��<@��<��<��<4��<r��<4��<	��<��<H��<\��<D��<@��<W��<e��<���<S��<r��<S��<���<e��<O��<@��<`   `   R��<h��<D��<P��<b��<N��<V��<k��<L��<>��<f��<R��<@��<I��<]��<K��<��<Z��<K��<��<W��<j��<D��<8��<`   `   5��<i��<C��<b��<&��<��<��<b��<N��<i��<5��<o��<W��<]��<���<���<?��<Q��<^��<���<j��<]��<d��<o��<`   `   W��<K��<?��<"��<!��<*��<*��<9��<G��<W��<?��<v��<e��<K��<���<؉�<[��<K��<ɉ�<���<W��<^��<p��<A��<`   `   ]��<9��<���<E��<W��<E��<���<9��<a��<F��<=��<Z��<���<��<?��<[��<\��<[��<A��<��<���<Z��<A��<F��<`   `   C��<P��<Z��<_��<V��<T��<Y��<D��<S��<U��<J��<E��<S��<Z��<Q��<K��<[��<^��<K��<K��<P��<L��<P��<W��<`   `   Z��<]��</��<S��<>��<]��<Q��<E��<6��<���<a��<���<r��<K��<^��<ɉ�<A��<K��<���<���<T��<���<7��<E��<`   `   U��<9��<F��<@��<1��<V��<R��<#��<o��<U��<T��<���<S��<��<���<���<��<K��<���<V��<`��<s��<��<J��<`   `   G��<?��<���<?��<O��<s��<e��<F��<���<`��<F��<P��<���<W��<j��<W��<���<P��<T��<`��<u��<F��<s��<s��<`   `   m��<K��<Q��<n��<l��<H��<m��<;��<o��<���<J��<K��<e��<j��<]��<^��<Z��<L��<���<s��<F��<e��<B��<u��<`   `   ��<	��<��<a��<
��<B��<v��<��<,��<P��<R��<p��<O��<D��<d��<p��<A��<P��<7��<��<s��<B��<��<a��<`   `   O��<P��<���<g��<l��<h��<R��<T��<S��<7��<?��<|��<@��<8��<o��<A��<F��<W��<E��<J��<s��<u��<a��<��<`   `   ��<���<��<���<���<���<���<���<���<���<���<���<ʈ�<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<��<���<���<ۈ�<���<���<���<���<҈�<È�<���<���<ň�<Ȉ�<���<���<���<���<߈�<���<���<
��<���<`   `   ��<���<���<ň�<���<���<ވ�<���<���<���<ψ�<���<ň�<���<���<���<ֈ�<���<���<ň�<���<���<���<���<`   `   ���<���<ň�<���<È�<���<���<ň�<���<È�<���<���<ʈ�<���<���<���<���<ǈ�<���<È�<���<���<߈�<��<`   `   ���<ۈ�<���<È�<݈�<ǈ�<���<��<݈�<���<���<���<Ո�<��<Ɉ�<ǈ�<͈�<È�<���<ۈ�<���<p��<���<p��<`   `   ���<���<���<���<ǈ�<���<���<���<���<���<���<���<���<���<��<ˈ�<���<���<���<���<���<ƈ�<���<���<`   `   ���<���<ވ�<���<���<���<���<���<���<���<���<���<���<���<�<���<Ԉ�<���<���<���<���<���<���<���<`   `   ���<���<���<ň�<��<���<���<߈�<ш�<҈�<݈�<���<���<��<���<���<���<���<���<���<���<|��<���<Ȉ�<`   `   ���<���<���<���<݈�<���<���<ш�<��<ш�<���<���<҈�<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<҈�<���<È�<���<���<���<҈�<ш�<���<���<ň�<ʈ�<���<Ȉ�<���<���<���<Ȉ�<t��<}��<ӈ�<���<���<`   `   ���<È�<ψ�<���<���<���<���<݈�<���<���<���<���<ʈ�<È�<���<���<���<t��<���<���<���<t��<���<���<`   `   ���<���<���<���<���<���<���<���<���<ň�<���<���<���<���<���<҈�<x��<���<���<���<���<m��<͈�<���<`   `   ʈ�<���<ň�<ʈ�<Ո�<���<���<���<҈�<ʈ�<ʈ�<���<ň�<���<���<���<ۈ�<���<T��<���<ވ�<���<���<���<`   `   ���<ň�<���<���<��<���<���<��<���<���<È�<���<���<���<���<���<���<ӈ�<Ȉ�<���<���<���<���<���<`   `   ���<Ȉ�<���<���<Ɉ�<��<�<���<���<Ȉ�<���<���<���<���<���<���<m��<ˈ�<���<���<���<���<���<���<`   `   ���<���<���<���<ǈ�<ˈ�<���<���<���<���<���<҈�<���<���<���<b��<���<���<V��<���<���<���<͈�<���<`   `   ���<���<ֈ�<���<͈�<���<Ԉ�<���<���<���<���<x��<ۈ�<���<m��<���<��<���<n��<���<و�<x��<���<���<`   `   ���<���<���<ǈ�<È�<���<���<���<���<���<t��<���<���<ӈ�<ˈ�<���<���<Ո�<Ȉ�<���<���<v��<���<���<`   `   ���<���<���<���<���<���<���<���<���<Ȉ�<���<���<T��<Ȉ�<���<V��<n��<Ȉ�<f��<���<���<Ȉ�<���<���<`   `   ���<߈�<ň�<È�<ۈ�<���<���<���<���<t��<���<���<���<���<���<���<���<���<���<���<}��<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<}��<���<���<ވ�<���<���<���<و�<���<���<}��<���<���<���<���<`   `   ���<���<���<���<p��<ƈ�<���<|��<���<ӈ�<t��<m��<���<���<���<���<x��<v��<Ȉ�<���<���<���<���<t��<`   `   ���<
��<���<߈�<���<���<���<���<���<���<���<͈�<���<���<���<͈�<���<���<���<���<���<���<���<߈�<`   `   ���<���<���<��<p��<���<���<Ȉ�<���<���<���<���<���<���<���<���<���<���<���<���<���<t��<߈�<���<`   `   L��</��<��<)��<X��<��<!��<C��<.��<(��<:��<@��<r��<@��<=��<(��<)��<C��<'��<��<S��<)��<��</��<`   `   /��<D��<��<B��<6��<9��<��<���<#��<2��<��<��<��<��<,��<!��< ��<��<3��<5��<H��<��<?��<,��<`   `   ��<��<%��<��<3��<J��<��<A��<��<��<6��</��<.��<��<#��<A��<��<J��<;��<��<��<��<��<Ї�<`   `   )��<B��<��<)��<3��<��<@��<1��<��<B��</��<2��<G��<��<+��<A��<
��<2��<"��<��<H��<&��<���<��<`   `   X��<6��<3��<3��<��<B��<��<��<*��<��<��<��<'��<��<��<B��<���<3��<8��<6��<U��<<��<Z��<<��<`   `   ��<9��<J��<��<B��<+��<��<4��<��<<��<9��<��<9��<��<%��<A��<
��<K��<3��<��<��<O��<K��<��<`   `   !��<��<��<@��<��<��<]��<5��<��<>��<��<5��<X��<��<	��<@��<��<��<+��<!��<��<���<��<!��<`   `   C��<���<A��<1��<��<4��<5��<��<��<��<��<6��<9��<��<+��<C��< ��<@��<9��<N��<X��<R��<J��<?��<`   `   .��<#��<��<��<*��<��<��<��<��<��<��<��<&��<��< ��<#��<*��<$��<��<6��<w��<6��<��<$��<`   `   (��<2��<��<B��<��<<��<>��<��<��<?��<9��<��<G��<��<,��<&��<"��<3��< ��<#��<)��<��</��<��<`   `   :��<��<6��</��<��<9��<��<��<��<9��<��</��<0��<��<C��<&��<Q��<i��<`��<���<S��<i��<\��<&��<`   `   @��<��</��<2��<��<��<5��<6��<��<��</��<1��<��<>��<��<��<9��<O��<>��<E��<U��<2��<��<!��<`   `   r��<��<.��<G��<'��<9��<X��<9��<&��<G��<0��<��<p��<&��<��<��<?��<-��<��<-��<@��<��<��<&��<`   `   @��<��<��<��<��<��<��<��<��<��<��<>��<&��<Q��<c��<��<:��<K��<E��<3��<��<i��<L��<!��<`   `   =��<,��<#��<+��<��<%��<	��<+��< ��<,��<C��<��<��<c��<J��<Q��<:��<F��<G��<Q��<>��<c��<'��<��<`   `   (��<!��<A��<A��<B��<A��<@��<C��<#��<&��<&��<��<��<��<Q��<X��<-��<'��<Q��<W��<��<��<��<)��<`   `   )��< ��<��<
��<���<
��<��< ��<*��<"��<Q��<9��<?��<:��<:��<-��<L��<-��<:��<:��<>��<9��<R��<"��<`   `   C��<��<J��<2��<3��<K��<��<@��<$��<3��<i��<O��<-��<K��<F��<'��<-��<L��<E��<(��<U��<l��</��<"��<`   `   '��<3��<;��<"��<8��<3��<+��<9��<��< ��<`��<>��<��<E��<G��<Q��<:��<E��<��<>��<W��< ��<��<9��<`   `   ��<5��<��<��<6��<��<!��<N��<6��<#��<���<E��<-��<3��<Q��<W��<:��<(��<>��<���<)��<4��<J��<"��<`   `   S��<H��<��<H��<U��<��<��<X��<w��<)��<S��<U��<@��<��<>��<��<>��<U��<W��<)��<s��<X��<��<��<`   `   )��<��<��<&��<<��<O��<���<R��<6��<��<i��<2��<��<i��<c��<��<9��<l��< ��<4��<X��< ��<K��<;��<`   `   ��<?��<��<���<Z��<K��<��<J��<��</��<\��<��<��<L��<'��<��<R��</��<��<J��<��<K��<_��<���<`   `   /��<,��<Ї�<��<<��<��<!��<?��<$��<��<&��<!��<&��<!��<��<)��<"��<"��<9��<"��<��<;��<���<҇�<`   `   ��<���<���<Շ�<���<���<���<Ň�<ڇ�<���<Շ�<���<���<���<Ӈ�<���<އ�<Ň�<���<���<���<Շ�<���<���<`   `   ���<f��<Ƈ�<���<V��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<Q��<���<ˇ�<d��<���<`   `   ���<Ƈ�<��<���<���<և�<���<���<͇�<���<���<ɇ�<���<���<Ӈ�<���<���<և�<���<���<އ�<Ƈ�<���<��<`   `   Շ�<���<���<���<���<�<Ç�<̇�<͇�<���<���<���<���<ȇ�<ˇ�<ȇ�<Ç�<���<���<���<���<ч�<݇�<߇�<`   `   ���<V��<���<���<���<���<���<ɇ�<���<���<χ�<���<���<ɇ�<���<���<���<���<���<V��<���<���<���<���<`   `   ���<���<և�<�<���<���<��<Ň�<���<݇�<ڇ�<���<Ǉ�<��<���<���<Ç�<ۇ�<���<���<Ň�<���<���<Ç�<`   `   ���<���<���<Ç�<���<��<���<���<���<���<���<���<���<��<���<Ç�<���<���<���<���<���<���<���<���<`   `   Ň�<���<���<̇�<ɇ�<Ň�<���<��<ʇ�<Ƈ�<���<���<Ǉ�<ć�<ˇ�<���<���<���<���<���<���<���<���<���<`   `   ڇ�<���<͇�<͇�<���<���<���<ʇ�<݇�<ʇ�<���<���<���<͇�<ʇ�<���<݇�<Ç�<���<���<���<���<���<Ç�<`   `   ���<���<���<���<���<݇�<���<Ƈ�<ʇ�<���<ڇ�<���<���<���<���<���<���<ć�<���<���<���<���<���<���<`   `   Շ�<���<���<���<χ�<ڇ�<���<���<���<ڇ�<ׇ�<���<���<���<ڇ�<���<���<���<q��<���<o��<���<���<���<`   `   ���<���<ɇ�<���<���<���<���<���<���<���<���<·�<���<���<ȇ�<���<���<h��<���<���<j��<���<���<ʇ�<`   `   ���<���<���<���<���<Ǉ�<���<Ǉ�<���<���<���<���<���<���<���<ڇ�<���<���<���<���<���<ڇ�<���<���<`   `   ���<���<���<ȇ�<ɇ�<��<��<ć�<͇�<���<���<���<���<���<���<���<���<���<���<���<���<���<��<}��<`   `   Ӈ�<���<Ӈ�<ˇ�<���<���<���<ˇ�<ʇ�<���<ڇ�<ȇ�<���<���<s��<���<���<q��<���<���<p��<���<���<ȇ�<`   `   ���<���<���<ȇ�<���<���<Ç�<���<���<���<���<���<ڇ�<���<���<߇�<���<���<އ�<���<���<ׇ�<���<���<`   `   އ�<���<���<Ç�<���<Ç�<���<���<݇�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   Ň�<���<և�<���<���<ۇ�<���<���<Ç�<ć�<���<h��<���<���<q��<���<���<s��<���<���<j��<���<���<���<`   `   ���<���<���<���<���<���<���<���<���<���<q��<���<���<���<���<އ�<���<���<���<���<l��<���<���<���<`   `   ���<Q��<���<���<V��<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<އ�<���<���<Ň�<���<���<���<���<o��<j��<���<���<p��<���<���<j��<l��<���<���<���<���<Ň�<`   `   Շ�<ˇ�<Ƈ�<ч�<���<���<���<���<���<���<���<���<ڇ�<���<���<ׇ�<���<���<���<���<���<���<���<���<`   `   ���<d��<���<݇�<���<���<���<���<���<���<���<���<���<��<���<���<���<���<���<���<���<���<���<݇�<`   `   ���<���<��<߇�<���<Ç�<���<���<Ç�<���<���<ʇ�<���<}��<ȇ�<���<���<���<���<���<Ň�<���<݇�<��<`   `   ��<$��<Y��<0��<Z��<���<C��<,��<M��<G��<5��<2��<j��<2��<.��<H��<X��<,��<6��<���<f��<0��<S��<$��<`   `   $��<`��<N��<5��<~��<V��<E��<o��<8��<2��<^��<g��<g��<a��<6��<2��<j��<M��<Z��<u��<2��<U��<`��< ��<`   `   Y��<N��<,��<���<K��<��<>��<8��<3��<j��<S��<Q��<Q��<j��<6��<8��<:��<��<N��<���<'��<N��<^��<Y��<`   `   0��<5��<���<\��<*��<k��<B��<��<7��<:��<9��<<��<:��<0��<��<J��<f��<"��<a��<���<2��<,��<B��<B��<`   `   Z��<~��<K��<*��<���<N��<K��<>��<Z��<R��<P��<R��<a��<>��<?��<N��<���<*��<?��<~��<a��<'��<6��<'��<`   `   ���<V��<��<k��<N��<I��<J��<0��<c��<-��<*��<\��<0��<S��<M��<E��<f��<$��<Z��<~��<A��<c��<c��<C��<`   `   C��<E��<>��<B��<K��<J��<��<K��<G��< ��<P��<K��<���<J��<P��<B��<<��<E��<C��<F��<X��<���<V��<F��<`   `   ,��<o��<8��<��<>��<0��<K��<���<4��<.��<���<T��<0��<5��<��<?��<j��<(��<=��<X��<L��<O��<W��<8��<`   `   M��<8��<3��<7��<Z��<c��<G��<4��<9��<4��<A��<c��<c��<7��<(��<8��<V��<4��<j��<F��<@��<F��<p��<4��<`   `   H��<2��<j��<:��<R��<-��< ��<.��<4��<	��<*��<I��<:��<r��<6��<C��<Z��<L��<g��<���<���<b��<L��<_��<`   `   5��<^��<S��<9��<P��<*��<P��<���<A��<*��<\��<9��<M��<^��<5��<r��<V��<g��<k��<`��<s��<g��<Q��<r��<`   `   2��<g��<Q��<<��<R��<\��<K��<T��<c��<I��<9��<X��<g��<.��<?��<N��<V��<u��<T��<O��<r��<[��<M��<;��<`   `   j��<g��<Q��<:��<a��<0��<���<0��<c��<:��<M��<g��<o��<���<P��<C��<d��<[��<Y��<[��<a��<C��<U��<���<`   `   2��<a��<j��<0��<>��<S��<J��<5��<7��<r��<^��<.��<���<}��<6��<���<q��<H��<L��<v��<���<2��<}��<���<`   `   .��<6��<6��<��<?��<M��<P��<��<(��<6��<5��<?��<P��<6��<i��<^��<g��<���<]��<^��<o��<6��<P��<?��<`   `   H��<2��<8��<J��<N��<E��<B��<?��<8��<C��<r��<N��<C��<���<^��<��<k��<p��<��<Z��<���<C��<M��<t��<`   `   X��<j��<:��<f��<���<f��<<��<j��<V��<Z��<V��<V��<d��<q��<g��<k��<C��<k��<f��<q��<f��<V��<T��<Z��<`   `   ,��<M��<��<"��<*��<$��<E��<(��<4��<L��<g��<u��<[��<H��<���<p��<k��<���<L��<\��<r��<j��<L��<.��<`   `   6��<Z��<N��<a��<?��<Z��<C��<=��<j��<g��<k��<T��<Y��<L��<]��<��<f��<L��<T��<T��<k��<g��<q��<=��<`   `   ���<u��<���<���<~��<~��<F��<X��<F��<���<`��<O��<[��<v��<^��<Z��<q��<\��<T��<c��<���<@��<W��<N��<`   `   f��<2��<'��<2��<a��<A��<X��<L��<@��<���<s��<r��<a��<���<o��<���<f��<r��<k��<���<I��<L��<P��<A��<`   `   0��<U��<N��<,��<'��<c��<���<O��<F��<b��<g��<[��<C��<2��<6��<C��<V��<j��<g��<@��<L��<���<c��<��<`   `   S��<`��<^��<B��<6��<c��<V��<W��<p��<L��<Q��<M��<U��<}��<P��<M��<T��<L��<q��<W��<P��<c��<?��<B��<`   `   $��< ��<Y��<B��<'��<C��<F��<8��<4��<_��<r��<;��<���<���<?��<t��<Z��<.��<=��<N��<A��<��<B��<`��<`   `   O��<(��<ۆ�<���<��<���<��<��<׆�<��<��<��<ӆ�<��<���<��<��<��<���<���<(��<���<ц�<(��<`   `   (��<+��<��<��<��<Ն�<��<��<	��<���<��<��<���<��<���<��<��<'��<߆�<��<	��<��<-��<#��<`   `   ۆ�<��<���<ц�<��<	��<��< ��<#��<���<ن�<��<ۆ�<���<"��< ��<��<	��<	��<ц�<���<��<ކ�<ֆ�<`   `   ���<��<ц�<ӆ�<��<��<	��<��<���<���<��<��<���<��<��<��<���<���<݆�<چ�<	��<���<��<��<`   `   ��<��<��<��<���<Ć�<)��<��<���<���<��<���<��<��<��<Ć�<��<��<��<��<!��<0��<W��<0��<`   `   ���<Ն�<	��<��<Ć�<��<��<��<���<���<���<��<	��<��<���<���<���<��<߆�<���<׆�<��<��<ކ�<`   `   ��<��<��<	��<)��<��<*��<1��<��<y��<���<1��<#��<��<,��<	��<��<��<��<���<���<͆�<���<���<`   `   ��<��< ��<��<��<��<1��<���<��<���<���<<��<	��<��<��<)��<��<���<;��<���<��<��<��<0��<`   `   ׆�<	��<#��<���<���<���<��<��<(��<��<��<���<��<���<��<	��<��<��<��<̆�<��<̆�<
��<��<`   `   ��<���<���<���<���<���<y��<���<��<���<���<��<���<��<���< ��<��<҆�<���<��<ކ�<���<ӆ�<��<`   `   ��<��<ن�<��<��<���<���<���<��<���<��<��<Ԇ�<��<��<��<���<��<��<ʆ�<���<��<��<��<`   `   ��<��<��<��<���<��<1��<<��<���<��<��<��<���<��<چ�<��<���<��<��<��<��<��<���<ц�<`   `   ӆ�<���<ۆ�<���<��<	��<#��<	��<��<���<Ԇ�<���<ۆ�<��<��<ن�<���<׆�<��<׆�<���<ن�<��<��<`   `   ��<��<���<��<��<��<��<��<���<��<��<��<��<���<���<���<���<Æ�<Ά�<���<��<��<���<��<`   `   ���<���<"��<��<��<���<,��<��<��<���<��<چ�<��<���<��<��<��<��<���<��<��<���<��<چ�<`   `   ��<��< ��<��<Ć�<���<	��<)��<	��< ��<��<��<ن�<���<��<���<��<��<Æ�<��<��<݆�<���<��<`   `   ��<��<��<���<��<���<��<��<��<��<���<���<���<���<��<��<Ć�<��<��<���<���<���<��<��<`   `   ��<'��<	��<���<��<��<��<���<��<҆�<��<��<׆�<Æ�<��<��<��<��<Ά�<چ�<��<��<ӆ�<��<`   `   ���<߆�<	��<݆�<��<߆�<��<;��<��<���<��<��<��<Ά�<���<Æ�<��<Ά�<׆�<��<��<���<��<;��<`   `   ���<��<ц�<چ�<��<���<���<���<̆�<��<ʆ�<��<׆�<���<��<��<���<چ�<��<̆�<ކ�<Ć�<��<��<`   `   (��<	��<���<	��<!��<׆�<���<��<��<ކ�<���<��<���<��<��<��<���<��<��<ކ�<&��<��<���<׆�<`   `   ���<��<��<���<0��<��<͆�<��<̆�<���<��<��<ن�<��<���<݆�<���<��<���<Ć�<��<؆�<��<$��<`   `   ц�<-��<ކ�<��<W��<��<���<��<
��<ӆ�<��<���<��<���<��<���<��<ӆ�<��<��<���<��<a��<��<`   `   (��<#��<ֆ�<��<0��<ކ�<���<0��<��<��<��<ц�<��<��<چ�<��<��<��<;��<��<׆�<$��<��<߆�<`   `   f��<���<���<���<���<���<ӆ�<���<���<���<ֆ�<��<���<��<ǆ�<���<Ɔ�<���<���<���<���<���<���<���<`   `   ���<e��<̆�<��<���<���<̆�<���<���<���<���<ц�<ʆ�<���<���<���<���<ن�<���<���<��<ֆ�<i��<���<`   `   ���<̆�<Ć�<׆�<���<҆�<b��<���<���<���<���<܆�<���<���<���<���<f��<҆�<���<׆�<ņ�<̆�<���<��<`   `   ���<��<׆�<���<���<׆�<���<���<���<ӆ�<Ά�<φ�<͆�<���<���<Ć�<ǆ�<���<���<��<��<���<�<���<`   `   ���<���<���<���<���<Ɔ�<���<���<ӆ�<���<���<���<��<���<Ɔ�<Ɔ�<φ�<���<߆�<���<���<���<���<���<`   `   ���<���<҆�<׆�<Ɔ�<���<���<���<���<���<���<���<���<���<Ɔ�<���<ǆ�<݆�<���<���<��<���<���<��<`   `   ӆ�<̆�<b��<���<���<���<���<Ȇ�<���<��<���<Ȇ�<���<���<��<���<h��<̆�<ǆ�<���<��<̆�<���<���<`   `   ���<���<���<���<���<���<Ȇ�<���<���<���<���<Ն�<���<���<���<���<���<���<~��<���<І�<ۆ�<���<n��<`   `   ���<���<���<���<ӆ�<���<���<���<ʆ�<���<���<���<��<���<���<���<�<���<��<���<���<���<��<���<`   `   ���<���<���<ӆ�<���<���<��<���<���<���<���<���<͆�<���<���<���<̆�<��<��<��<߆�<��<���<݆�<`   `   ֆ�<���<���<Ά�<���<���<���<���<���<���<���<Ά�<���<���<͆�<���<���<���<���<���<ۆ�<���<x��<���<`   `   ��<ц�<܆�<φ�<���<���<Ȇ�<Ն�<���<���<Ά�<��<ʆ�<��<Ն�<͆�<ކ�<���<���<���<���<��<ц�<Ȇ�<`   `   ���<ʆ�<���<͆�<��<���<���<���<��<͆�<���<ʆ�<���<�<܆�<	��<���<ކ�</��<ކ�<���<	��<��<�<`   `   ��<���<���<���<���<���<���<���<���<���<���<��<�<���<Ɔ�<ʆ�<��<̆�<ۆ�<���<���<���<���<Ɇ�<`   `   ǆ�<���<���<���<Ɔ�<Ɔ�<��<���<���<���<͆�<Ն�<܆�<Ɔ�<���<���<��<d��<҆�<���<���<Ɔ�<ц�<Ն�<`   `   ���<���<���<Ć�<Ɔ�<���<���<���<���<���<���<͆�<	��<ʆ�<���<��<؆�<��<��<���<���<��<ц�<���<`   `   Ɔ�<���<f��<ǆ�<φ�<ǆ�<h��<���<�<̆�<���<ކ�<���<��<��<؆�<ˆ�<؆�<���<��<���<ކ�<���<̆�<`   `   ���<ن�<҆�<���<���<݆�<̆�<���<���<��<���<���<ކ�<̆�<d��<��<؆�<W��<ۆ�<��<���<���<���<���<`   `   ���<���<���<���<߆�<���<ǆ�<~��<��<��<���<���</��<ۆ�<҆�<��<���<ۆ�<��<���<ˆ�<��<��<~��<`   `   ���<���<׆�<��<���<���<���<���<���<��<���<���<ކ�<���<���<���<��<��<���<���<߆�<���<���<��<`   `   ���<��<ņ�<��<���<��<��<І�<���<߆�<ۆ�<���<���<���<���<���<���<���<ˆ�<߆�<Ɇ�<І�<ކ�<��<`   `   ���<ֆ�<̆�<���<���<���<̆�<ۆ�<���<��<���<��<	��<���<Ɔ�<��<ކ�<���<��<���<І�<ن�<���<���<`   `   ���<i��<���<�<���<���<���<���<��<���<x��<ц�<��<���<ц�<ц�<���<���<��<���<ކ�<���<���<�<`   `   ���<���<��<���<���<��<���<n��<���<݆�<���<Ȇ�<�<Ɇ�<Ն�<���<̆�<���<~��<��<��<���<�<)��<`   `   چ�<���<���<���<x��<���<���<���<���<���<���<d��<O��<d��<���<���<���<���<���<���<���<���<���<���<`   `   ���<���<���<���<���<h��<���<ن�<���<|��<���<���<}��<���<���<���<Ć�<���<|��<���<���<���<���<���<`   `   ���<���<��<���<���<i��<l��<���<ņ�<���<{��<���<���<���<���<���<r��<i��<���<���<��<���<���<���<`   `   ���<���<���<Y��<W��<φ�<���<X��<���<���<\��<\��<w��<��<i��<ˆ�<���<H��<m��<���<���<���<���<~��<`   `   x��<���<���<W��<���<q��<���<���<���<���<���<���<���<���<x��<q��<���<W��<���<���<���<|��<���<|��<`   `   ���<h��<i��<φ�<q��<R��<Ć�<���<���<���<���<���<���<ӆ�<b��<b��<���<u��<|��<���<���<���<���<���<`   `   ���<���<l��<���<���<Ć�<L��<���<���<J��<���<���<G��<Ć�<���<���<u��<���<���<���<m��<���<Y��<���<`   `   ���<ن�<���<X��<���<���<���<���<���<w��<���<���<���<��<i��<ņ�<Ć�<���<\��<f��<���<���<l��<H��<`   `   ���<���<ņ�<���<���<���<���<���<���<���<���<���<���<���<���<���<���<t��<���<���<6��<���<���<t��<`   `   ���<|��<���<���<���<���<J��<w��<���<X��<���<w��<w��<Æ�<���<���<���<Z��<f��<���<y��<R��<`��<���<`   `   ���<���<{��<\��<���<���<���<���<���<���<���<\��<y��<���<���<���<���<e��<x��<���<���<e��<k��<���<`   `   d��<���<���<\��<���<���<���<���<���<w��<\��<���<}��<a��<p��<e��<���<���<`��<M��<���<Æ�<j��<_��<`   `   O��<}��<���<w��<���<���<G��<���<���<w��<y��<}��<[��<���<]��<^��<Q��<c��<n��<c��<K��<^��<h��<���<`   `   d��<���<���<��<���<ӆ�<Ć�<��<���<Æ�<���<a��<���<���<z��<���<���<P��<d��<���<���<i��<���<���<`   `   ���<���<���<i��<x��<b��<���<i��<���<���<���<p��<]��<z��<���<i��<���<m��<y��<i��<چ�<z��<N��<p��<`   `   ���<���<���<ˆ�<q��<b��<���<ņ�<���<���<���<e��<^��<���<i��<O��<���<���<c��<X��<���<g��<j��<���<`   `   ���<Ć�<r��<���<���<���<u��<Ć�<���<���<���<���<Q��<���<���<���<%��<���<���<���<V��<���<��<���<`   `   ���<���<i��<H��<W��<u��<���<���<t��<Z��<e��<���<c��<P��<m��<���<���<\��<d��<l��<���<f��<`��<k��<`   `   ���<|��<���<m��<���<|��<���<\��<���<f��<x��<`��<n��<d��<y��<c��<���<d��<R��<`��<���<f��<���<\��<`   `   ���<���<���<���<���<���<���<f��<���<���<���<M��<c��<���<i��<X��<���<l��<`��<���<y��<y��<l��<���<`   `   ���<���<��<���<���<���<m��<���<6��<y��<���<���<K��<���<چ�<���<V��<���<���<y��<M��<���<Y��<���<`   `   ���<���<���<���<|��<���<���<���<���<R��<e��<Æ�<^��<i��<z��<g��<���<f��<f��<y��<���<���<���<m��<`   `   ���<���<���<���<���<���<Y��<l��<���<`��<k��<j��<h��<���<N��<j��<��<`��<���<l��<Y��<���<Ć�<���<`   `   ���<���<���<~��<|��<���<���<H��<t��<���<���<_��<���<���<p��<���<���<k��<\��<���<���<m��<���<���<`   `   ���<L��<a��<���<u��<k��<���<q��<��<V��<���<h��<h��<h��<���<V��<=��<q��<j��<k��<���<���<N��<L��<`   `   L��<p��<���<���<c��<5��<b��<t��<)��<@��<u��<���<���<u��<S��< ��<]��<r��<K��<R��<���<���<v��<I��<`   `   a��<���<=��<���<���<���<��<p��<���<���<c��<���<m��<���<w��<p��<��<���<���<���<B��<���<]��<��<`   `   ���<���<���<i��<���<���<x��<M��<T��<���<|��<|��<u��<K��<`��<���<���<|��<���<���<���<���<_��<X��<`   `   u��<c��<���<���<o��<M��<���<f��<R��<O��<���<O��<f��<f��<o��<M��<���<���<���<c��<���<v��<�<v��<`   `   k��<5��<���<���<M��<>��<���<���<J��<z��<{��<A��<v��<���<Q��<=��<���<���<K��<g��<[��<e��<l��<k��<`   `   ���<b��<��<x��<���<���<,��<>��<R��<j��<[��<>��<'��<���<���<x��<!��<b��<|��<v��<;��<r��<#��<v��<`   `   q��<t��<p��<M��<f��<���<>��<Q��<m��<d��<Q��<M��<v��<V��<`��<{��<]��<n��<���<���<���<���<���<���<`   `   ��<)��<���<T��<R��<J��<R��<m��<ņ�<m��<C��<J��<m��<T��<b��<)��<7��<m��<Ć�<���<i��<���<Ԇ�<m��<`   `   V��<@��<���<���<O��<z��<j��<d��<m��<z��<{��<?��<u��<���<S��<S��<~��<S��<@��<���<���<)��<Z��<���<`   `   ���<u��<c��<|��<���<{��<[��<Q��<C��<{��<���<|��<a��<u��<���<���<���<���<p��<���<���<���<r��<���<`   `   h��<���<���<|��<O��<A��<>��<M��<J��<?��<|��<���<���<e��<g��<v��<���<���<~��<h��<���<���<}��<T��<`   `   h��<���<m��<u��<f��<v��<'��<v��<m��<u��<a��<���<v��<���<���<o��<>��<���<ņ�<���<7��<o��<���<���<`   `   h��<u��<���<K��<f��<���<���<V��<T��<���<u��<e��<���<���<c��<���<���<c��<z��<���<���<O��<���<���<`   `   ���<S��<w��<`��<o��<Q��<���<`��<b��<S��<���<g��<���<c��<���<c��<���<���<w��<c��<���<c��<���<g��<`   `   V��< ��<p��<���<M��<=��<x��<{��<)��<S��<���<v��<o��<���<c��<7��<���<���<N��<P��<���<y��<}��<���<`   `   =��<]��<��<���<���<���<!��<]��<7��<~��<���<���<>��<���<���<���<��<���<���<���<D��<���<���<~��<`   `   q��<r��<���<|��<���<���<b��<n��<m��<S��<���<���<���<c��<���<���<���<���<z��<���<���<���<Z��<c��<`   `   j��<K��<���<���<���<K��<|��<���<Ć�<@��<p��<~��<ņ�<z��<w��<N��<���<z��<���<~��<���<@��<ǆ�<���<`   `   k��<R��<���<���<c��<g��<v��<���<���<���<���<h��<���<���<c��<P��<���<���<~��<���<���<���<���<���<`   `   ���<���<B��<���<���<[��<;��<���<i��<���<���<���<7��<���<���<���<D��<���<���<���<���<���<$��<[��<`   `   ���<���<���<���<v��<e��<r��<���<���<)��<���<���<o��<O��<c��<y��<���<���<@��<���<���<���<l��<f��<`   `   N��<v��<]��<_��<�<l��<#��<���<Ԇ�<Z��<r��<}��<���<���<���<}��<���<Z��<ǆ�<���<$��<l��<ˆ�<_��<`   `   L��<I��<��<X��<v��<k��<v��<���<m��<���<���<T��<���<���<g��<���<~��<c��<���<���<[��<f��<_��<$��<`   